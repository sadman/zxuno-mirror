-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0C330C320081FFFFD43FF5684402617B44017FFFFFFFFFFFF9FFFB120A301015";
    attribute INIT_01 of inst : label is "6152175124A81FA89A0049202900BEFE530D98942FA12A51FFFFFFFC6019009B";
    attribute INIT_02 of inst : label is "C41549F4FE1149F79E11E4C6989312624C7EEE016110B1A80322C50A16DFB9EE";
    attribute INIT_03 of inst : label is "24443C0500F0F6B4FB322A10D69F6654421A93ECC01843527D984328A02AF7D4";
    attribute INIT_04 of inst : label is "E7C185123F280087CDF4DC229442A9504FCA00214F054873C1523C050087CA02";
    attribute INIT_05 of inst : label is "00451555A856A15A8B6B84617A4A051738FFF9FFE75CF9337FC994067C185122";
    attribute INIT_06 of inst : label is "9201095010500800045554245490084A828A904008A2AAA122A4804254145482";
    attribute INIT_07 of inst : label is "1149420002D000B4004141114AF91108F8A4E08A1842AA86062AA1800AAA848A";
    attribute INIT_08 of inst : label is "154428ACBBD413012A022344A38B80010A11554BFC43FC0AA088008508A2B095";
    attribute INIT_09 of inst : label is "97D51C44F89FA3A0297F4739141FE2910B1AC6B0820495E4DB3D4138B8212881";
    attribute INIT_0A of inst : label is "6DB6C4D0C6DCDB1B6370FF47FA83FC5BF9DD22EE9577403BA11F3A2FF0060413";
    attribute INIT_0B of inst : label is "8FC42AA710AE1C42A8F12AE3CC1CFB72E5CDC18B163702A62C58DC18B1637008";
    attribute INIT_0C of inst : label is "5438207882FF7B1A3F7B39A300731981400AF576AB530431410D44800FE2A22A";
    attribute INIT_0D of inst : label is "77FFEC2DFA8840A5FD1EAF78D45054E87FB0B7E010007616F78040009D85B125";
    attribute INIT_0E of inst : label is "BFC4D47FA0FF4294ED6666666666666666666666666666A60CF9F3E73E7D85BF";
    attribute INIT_0F of inst : label is "49C6A1221FF081F3C93AA1236E468E83F2360280A44C1BFF3DFB88CE66CE5FB4";
    attribute INIT_10 of inst : label is "51DCFF7FD651328C2222424820A1010A05250000044812810848128108481281";
    attribute INIT_11 of inst : label is "D5B2F08409CFA2113A98000ACE74EF48EA2131CCDCED25E473FFDAE8AA84ACE7";
    attribute INIT_12 of inst : label is "FF201864E4A80224500844029A2A405429A4A69782A768BCE55466963695488C";
    attribute INIT_13 of inst : label is "D80C1A1185F1029228127962004A3A73E47E87CEE00000017FB78F1772577BDE";
    attribute INIT_14 of inst : label is "33CDFD05D73001DB2E187A0FBC5501401500A4950088878289A1183603068460";
    attribute INIT_15 of inst : label is "9BFDC877FD840352E7B17735763DEDEF7F9A08000017952119D5C08C83D7D5A6";
    attribute INIT_16 of inst : label is "555515528A850DA1554000E3598AA29C0AE24538B9516BA52F04458AB2A8B1A7";
    attribute INIT_17 of inst : label is "D215856058160585434090350D4258D4343BDB93FF308650444D6A110B36A855";
    attribute INIT_18 of inst : label is "AC5FF323FFFFF5DFFFFFFE0000000031A000096000BD278126266027299AD960";
    attribute INIT_19 of inst : label is "E621CBFB10E4FCDFD4FC3CCD49CDC026C799EDCF1040900E5C2103E4F73C9BFF";
    attribute INIT_1A of inst : label is "41FAC6F7B7C9BEE2054005E5F5F1F084BE11F10E5C5EEE0290026624912C4393";
    attribute INIT_1B of inst : label is "D8000008956DFEE915593EEFE977FEFFFFE96365D16087CBE5F2F97C87F43D0F";
    attribute INIT_1C of inst : label is "2222220200888880008888881BBFB7F75DB3970E9AE44F5DAC6DE6938047F745";
    attribute INIT_1D of inst : label is "0000000000000041000000000000088000028808880800008200008022222000";
    attribute INIT_1E of inst : label is "55555555555555555555555540400000020A08080C4500000000000000000041";
    attribute INIT_1F of inst : label is "7CDB379B4C6B75B212DE33BDEC952F3084046551451115150111111275757575";
    attribute INIT_20 of inst : label is "02A412D4884405373846B9EF6B3468E65CC19C7C8840A50A5CCF7F7DDFF7FDF7";
    attribute INIT_21 of inst : label is "F3FD3E2F801695A7C34A7C48D30F87C0AA7C3602040422452D30F86C0A53E1E4";
    attribute INIT_22 of inst : label is "05542FE9BD08D35845EB2383129B240F31ED9E23D09EFA4F5B3169259EC64431";
    attribute INIT_23 of inst : label is "FFB80FFFFF7FFFFFED878E01FE03FE03FF504E9D111111111111171C95AAB000";
    attribute INIT_24 of inst : label is "C716DF38A28A39F6F1C7CC79F5FFBC1EF9EEB7DAB7FFFFFEFF07FEFFFFFFC7FF";
    attribute INIT_25 of inst : label is "1F3DFFFFFF03BFEA03FFFF7BEFBBEDBEB3DF6CFB8E4BFFFBDFDBFEFAFF77EFF7";
    attribute INIT_26 of inst : label is "078E3FFCFB4D3FBC0F75FE7FDFFC7F47B7FFC7FFE57DE773070039E60E0073CF";
    attribute INIT_27 of inst : label is "7FFFFFFFF83F23F83F23F83F23F1FFFFFFFFFFFFFFFFFFF8F1FFF02F09F31C31";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "4D13423010A8FFFF0A404365B58F64F22244C03FFFFFFFFFF9FFEBF5318E7993";
    attribute INIT_01 of inst : label is "EDD81E5D86EC8AA40C4965B6EC927A6D18324B5E61370568FFFFFFF802184918";
    attribute INIT_02 of inst : label is "0A56140120522201205238CD19A334668CE61245E59BB6E65E26CD676A457FFE";
    attribute INIT_03 of inst : label is "B7DCE049900F0A5D181B30274BA3036600E9346064501D268C0C88233649D357";
    attribute INIT_04 of inst : label is "6012563B20B299C822284244212A4232782CA47200976CB0059BA04990DB6BB9";
    attribute INIT_05 of inst : label is "9167759CB972E5CB9D34972DA9670C880AFF0BFFBFAC0064FFD25924012563B3";
    attribute INIT_06 of inst : label is "DB24ECA134D962448DD6289092D927250BAED9122CE6914584B6C93B285D76D8";
    attribute INIT_07 of inst : label is "8C8488444BD948F65325C59929582020B2ECC9B33963AC4E486933921AC51612";
    attribute INIT_08 of inst : label is "8D75BCD0255D8D64B9491893A78F99132ED9D8AFFF67FF66724489976CCC625C";
    attribute INIT_09 of inst : label is "5D9DD8C844080A8CECD7280A5DFFE6DD94BFFF7279165C8052D5DCF8F997834C";
    attribute INIT_0A of inst : label is "4924A392AAD15A2B456D4D7FFBBFFC924AE5B372D9B9645CB22B233AA99D6970";
    attribute INIT_0B of inst : label is "523348B0CD22433C890CD22438A1A0448911B152A556E3B448911B1122456E19";
    attribute INIT_0C of inst : label is "D9082A0849C04102404120242618381322733DE8CDC8CC04949D23249AE6E6E6";
    attribute INIT_0D of inst : label is "93FE04A403ADD663C23110A3222627290412902C88C8825214B22322A094882C";
    attribute INIT_0E of inst : label is "FFF832FFE5FFCEE16C3333333333333333333333333333A3055A95687F009483";
    attribute INIT_0F of inst : label is "2D4096956AA3B1081403C2A4324AFF17F6444644F68138AA29526D2002E3DE3F";
    attribute INIT_10 of inst : label is "8A31044840C78639060D2B994532B4AF2893B6F24DED694A2CED694A6DAD694A";
    attribute INIT_11 of inst : label is "B880AB1D8463333692691966118A118B0EB77631023245F48C41192396326110";
    attribute INIT_12 of inst : label is "6C43422706ECCF9CDCF12231C66D7625917645C940035C429944B5C113048416";
    attribute INIT_13 of inst : label is "664DC4D9B263899914C88B06488BFC8AE9013C13000000013680182841584010";
    attribute INIT_14 of inst : label is "345A8B92CF2019080B000B1129A2928A4A29000601090205044D9B9BB371726E";
    attribute INIT_15 of inst : label is "648209843248CA058042840588610008320B550000101532814771D29ADB2175";
    attribute INIT_16 of inst : label is "666626622A8419328B000165806864A058D0C940346DA0469AB34D8E6A69B3FC";
    attribute INIT_17 of inst : label is "3DEA5B9FA5F9FA5B9CBD3FCA539CA579CA7C360C02C1F949CF724459242B3066";
    attribute INIT_18 of inst : label is "D08000DC00000A080000000000000000C00011200110AC0174046174C91B959D";
    attribute INIT_19 of inst : label is "456A2022B510123FDFFC9EE49A1C646AD3DCD5A6B52B5A511247621100C120C9";
    attribute INIT_1A of inst : label is "82A1207CC8160D07455004046E6A6E464DCA6B5110CD1D695A59927373EAD444";
    attribute INIT_1B of inst : label is "600000228049D904978320302AD8300C43108901488E64120904824105485214";
    attribute INIT_1C of inst : label is "7774754E5FDD1D5319DDD1D53284385120A86DC26486A444FAB09514A45116F4";
    attribute INIT_1D of inst : label is "BAAAAEBAEBAEBEAEBAAAAEBAEBAEB887D2249171D52859969F599797F74754C6";
    attribute INIT_1E of inst : label is "000000000202020200000000414000000008080838641088AA4222A9088AAEAE";
    attribute INIT_1F of inst : label is "0244C3400682012632A6000609064933C4004223A979797BA939393A00000000";
    attribute INIT_20 of inst : label is "DB369BA818D59D8685FDF3BDEF95DB80CF63DA25EDDA779685FE85024058040D";
    attribute INIT_21 of inst : label is "97FD94E5347B37529D9B29ABA934BA56EF29D2BB9859B369BA934BA56F794E8D";
    attribute INIT_22 of inst : label is "0554205FFA6CEB820F79CC953C4CCCB5DF79EBBEF1E097FE8CC7B336023708D6";
    attribute INIT_23 of inst : label is "11BAE00055D555001A9800000000000001B0850941414141414140A92701F000";
    attribute INIT_24 of inst : label is "00000000410400000001520609001BE10C1140049804000000F8000000400C10";
    attribute INIT_25 of inst : label is "106698003FFC456AA80A2816186413414C229B04308400040000040400000001";
    attribute INIT_26 of inst : label is "F05050036DB0D0BEF09A698004038838400838009B4001F0C00000018000000A";
    attribute INIT_27 of inst : label is "7FFFFFFFF83F03F83F03F83F03F1000000000000000000074E03FFF0F6082082";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "651943710DB8FFFF0202F1E02403414B54207FFFFFFFFFFFF8FFE06333045D01";
    attribute INIT_01 of inst : label is "40170641760C5C2B7A8201002000AFBB450DD8523EA5A14FFFFFFFFD21B8C0C8";
    attribute INIT_02 of inst : label is "421442442510504505102A8550AA1543A875D4A84C40F0A8C3AA85430DDA2508";
    attribute INIT_03 of inst : label is "B9C8DE458000001DB5188E5003B6A3114A0076D46229C00EDA8C4518240A6DD4";
    attribute INIT_04 of inst : label is "E2A09038950489C1FBEAEAABBD5ABA673541207107916271C4189E458A434BB3";
    attribute INIT_05 of inst : label is "99455527889EAA788B7D31C4710A15515AAA0F556DDD62756A9482182A09138C";
    attribute INIT_06 of inst : label is "02092121155A1A6514501C8C9082030908A2C0D3202282E564A0825A48455696";
    attribute INIT_07 of inst : label is "506516865082502094284C454A592120BE3AF8E0191820165688219182899192";
    attribute INIT_08 of inst : label is "41140E07B7D55D080AC88EDFAB6B50214244492AA94AA942922010A12224A005";
    attribute INIT_09 of inst : label is "D5D41D42E6EFE96021562D5A55354AD5A11294A4919040574BFD57F6B5219844";
    attribute INIT_0A of inst : label is "AEBAC2954EA9D53AB749534D52A6A94B5A09AA04D5026A81354BAAA559526F55";
    attribute INIT_0B of inst : label is "5F2243928B0E4A243B2890E4A935AFA74E9D2A9D3A64A28B76EDD2A9D3A64A28";
    attribute INIT_0C of inst : label is "DF0B6E0882E7D00A27D1482200FF1A8020145532A957C6FC3D2D56210ACE4646";
    attribute INIT_0D of inst : label is "935520A0C2A954A5F753A9C275F5F50804828328C8CC905072A32332B4140A68";
    attribute INIT_0E of inst : label is "2ABD60D541AA94306800F0F0F0F4F00F000F96FF0F0F0F0F05AB56AD75A41413";
    attribute INIT_0F of inst : label is "2086A08C655D169FDA50E5A82E529B0EA642AAEC7ED5515515ABCDE2A0028087";
    attribute INIT_10 of inst : label is "17D771058FB1FD8FEA095A9A4904AD2B4820841084694A52606108C221294AD2";
    attribute INIT_11 of inst : label is "7180A368B7D1AA548A82CA4BDEB0E32AEAA575C71C77D7E5758CAFE2A584BDEA";
    attribute INIT_12 of inst : label is "15F0FFF7F60C01FC541B1008FE29323434E6D39A80F639CC4429E38A77E1A2BC";
    attribute INIT_13 of inst : label is "A4E8748D0030C09885AEDA22624AF2892D1B85F7000000001B778F0F915791F4";
    attribute INIT_14 of inst : label is "96D12187142032180A082906B93284CA13282B03008C84850759D0F93A1F2743";
    attribute INIT_15 of inst : label is "EAFF6AD5E40A99D72BB0F915723F45F20CF87C000050052AE60F04C3B4AF8838";
    attribute INIT_16 of inst : label is "8787807888041AE28000014A85A589120821D224080D7F648F91514A320AA007";
    attribute INIT_17 of inst : label is "484291AD6B4A5291AD6B4A5295AD6B0A52A1C4CCB8991B44D087404149ABC07F";
    attribute INIT_18 of inst : label is "11ABF15C00000AA000000E000000005AC000088000A71E40330BC03222F1AA83";
    attribute INIT_19 of inst : label is "6253C2B129E15BBA85A821083B5AE214A4212D496918421E04DA2D3DF11D2B32";
    attribute INIT_1A of inst : label is "FB5AAA8519F6B223000414009692963612C6969E1552AA5A529E94BD7224A785";
    attribute INIT_1B of inst : label is "A800000A94422A64557F55FFCBCBD675DD758B01440D7BDDEEF77BBDFABF6FDB";
    attribute INIT_1C of inst : label is "7776770E5FDD9DC30DDDD9DC33D2AAFEDB3D7F9DB6F6EF7B5FD9F796402AB566";
    attribute INIT_1D of inst : label is "BAAAAAAAAAAAAEEFBAAAAAAAAAAAA897C5568D79DC2950C28750C397F76770C3";
    attribute INIT_1E of inst : label is "55555555575757575555555540400000000A0808286FEFAFFFBEBFFEFAFFFEEF";
    attribute INIT_1F of inst : label is "BF29D4AF50A8440732494107E94749024CAEC003EDB9BDBFA9B9B9BA75757575";
    attribute INIT_20 of inst : label is "4AA4CA0BA888016474562509426408AACAB3D5604956B4AF85B9783E0FCBF2F8";
    attribute INIT_21 of inst : label is "16A906A1A8583410D41A0D4A0850A954A90D4AA91454AA4CA0850A9549486A4D";
    attribute INIT_22 of inst : label is "80000755E5464D3BD5A86B17684368A2A9A94553534ED57943659394DF34C154";
    attribute INIT_23 of inst : label is "00B91000008000021DC00E01FE03FE03FE11C8900154015401540698F35CE000";
    attribute INIT_24 of inst : label is "8028004041044008028052060A0060000283005298007C0120FA01007C002690";
    attribute INIT_25 of inst : label is "004208003F00402A54000198000003800000000041240044202405150088100D";
    attribute INIT_26 of inst : label is "0082901B041240BD004105B8144041BC5BC104045A280D80C000000180000180";
    attribute INIT_27 of inst : label is "7FFFFFFC000000000000000002090020C00C0000040000064E03F0300004C34C";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "A29883585520FFFF8342B0C420E226791224543FFFFFFFFFF8FFF8299DEA0481";
    attribute INIT_01 of inst : label is "2423C48C256ADE475BB44800B0C22E9BCBA4F8422D812189FFFFFFFE0AA82CC0";
    attribute INIT_02 of inst : label is "4267425425A3505505A365ECAD953AE654E550246C4862865B04EA6F65B230AC";
    attribute INIT_03 of inst : label is "DEAEE56D5000010DF514D2B021BEA29A520437D4534AC086FA8A695880736CE2";
    attribute INIT_04 of inst : label is "C0AAAB75C55553AFEACAC227BD58FB2BB95556EBC15B556056D5C56D545E977F";
    attribute INIT_05 of inst : label is "158A20F9F7E7579D564942D09422484F5855C8FFC3591A21FFC6AAAA0AAAA754";
    attribute INIT_06 of inst : label is "F7DF2A34A3974C573987D8ACA73CFB51A51CBA62B9CC3CC4651965988D28A543";
    attribute INIT_07 of inst : label is "59E5D2EDFADE3A978E2D5D5C61B2EFEF5966659AD3DF4EA4E7538939D4791594";
    attribute INIT_08 of inst : label is "4C60AAFC95D9DD082A589AB51EECD8E2EAD58F7954795462962471756AC6B015";
    attribute INIT_09 of inst : label is "D6FECFEEE6EFEB68CD6CAF583D1FFCBD7FDC6717B7471F77595D9D6ECDA1384C";
    attribute INIT_0A of inst : label is "A69A536745E8AD97A2AD5F47FF23FF8959B96FDCB7EE5BF72DF61AB5595AAE55";
    attribute INIT_0B of inst : label is "5BA3AEF88CBB6232FF88CBF62D3CABA3468ABE8D1A2EFF5A3468ABECD9B2EFF5";
    attribute INIT_0C of inst : label is "B4114826689750C45710ACC584BF96C391606892250DE4DE516A773A4D9DFFDD";
    attribute INIT_0D of inst : label is "31FE6AE0222D16868F3399E1F676761111AB80821EE8B5701B087BA33D5C184A";
    attribute INIT_0E of inst : label is "3FE1402AC055843412F0FF00FF00FFF0000FFFFFF00FF00F09B3668F2BAD5C09";
    attribute INIT_0F of inst : label is "85AD18C7755CB89A98585147298E06A3F26224576ED41B55D4A945DAA21B0085";
    attribute INIT_10 of inst : label is "33C575C58AB5D5A8BA39CECB19A4E77BDF48E91D2579CE738579CEF384318CE3";
    attribute INIT_11 of inst : label is "3548BBE1C54489D0AC52AB035EA3E221E8B427D53D575358F14C8B4085A1B7EB";
    attribute INIT_12 of inst : label is "15BA6F77256AA9BD8A9B57AADEC7BAB98C663184001618682200A19001686114";
    attribute INIT_13 of inst : label is "ED4DDDA8B0945ABABCCAF8AF55F1CC410C879DD50000000059778F0F589F19C4";
    attribute INIT_14 of inst : label is "87C6B512045810500A8E39D29D2214895221A12A848883848D5A8BBB53776A2E";
    attribute INIT_15 of inst : label is "8A7C5355C75F0D763390F589F63C45E30AD8680000000131D6B0E59F153BA6AB";
    attribute INIT_16 of inst : label is "07F8007808115C22590001C0D402000A0803C014010A4D7485D31FEA1C635A97";
    attribute INIT_17 of inst : label is "BFEF7AD7B5ED7B5BFEF7FDFFFAD7B5EF6BCFD0AAFE546A0C9ABFC64861580078";
    attribute INIT_18 of inst : label is "99EB995C0000000000000E000000008180004A0004820E802101C0211071C0F7";
    attribute INIT_19 of inst : label is "FAD3C4F569E37EBFE8FEC5721BCAD35538AE2A71698C631E24F97135AD1F4D2A";
    attribute INIT_1A of inst : label is "C35F031671D2D332000000011717172B62E316BE2762D3CEF39A19B43CF4AF8D";
    attribute INIT_1B of inst : label is "A800000084002A64A7EE957E5353E4795E55CA9144E61BD9ECF67B3D82BC7F1F";
    attribute INIT_1C of inst : label is "2221201A088848064C88848079F8CB32491F93E4B26EF28946CE69A753BA28C2";
    attribute INIT_1D of inst : label is "504104545145151450410454514519D20771C424806D0CC3CA0CC28222120193";
    attribute INIT_1E of inst : label is "20202020020202022020202048CA0681A01DDF5D680BBB2200EC8803B2200514";
    attribute INIT_1F of inst : label is "BC2F14AD40884D0355575487080F0AB706104081135753511313171200000000";
    attribute INIT_20 of inst : label is "CABC2F0EE8898230D46291A4612088E2431527604973BCE4E445F43D0F0BC2F0";
    attribute INIT_21 of inst : label is "515586A1AF6C1610D60B0D7308DAAC46B90D6A3956DCABC2F08DAAD469C86B05";
    attribute INIT_22 of inst : label is "00000F07165C45EB74A86B162E416CBEACAE7559557E41C58167C1D6D6226F77";
    attribute INIT_23 of inst : label is "3F47F0000000000210000C01FE000000008C8000540001555400028C23906000";
    attribute INIT_24 of inst : label is "000000000100000000021206080000000082005200007C0000F800007C002210";
    attribute INIT_25 of inst : label is "0002080FC0FC0FD5FC0001800000038000000000002000000000041000000000";
    attribute INIT_26 of inst : label is "0000801B04107F43F04105B02000413C13C104045A280000C000000180000180";
    attribute INIT_27 of inst : label is "7FFFFFFC000000000000000002080000000C00000400000400FC0FF000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "340D0329D4E4FFFF6B52E2E4B4E404B07666957FFFFFFFFFF8FFE7AD11DA65AA";
    attribute INIT_01 of inst : label is "4494C94D5162E427216D6D9254D2D9449EB8235AD25AD52CFFFFFFFE7A902DEC";
    attribute INIT_02 of inst : label is "98D29809A0968A09A096448891502244488094ED85DB77244EA6093B7B200408";
    attribute INIT_03 of inst : label is "14CCC06850000559A105D082AB3420BA1455668417428AACD082E8515AC9DA16";
    attribute INIT_04 of inst : label is "6D1A4B25C8D2D928822B4265693253333234964AD89B15B626C5C0E85E4B5111";
    attribute INIT_05 of inst : label is "11AA6598FF63FD8FF0920601806CD9D95100A055406DAB04AA9269AAD1A5B255";
    attribute INIT_06 of inst : label is "FDF6ACB6AA8564C6A996B9BBD7EFB765B5542B22354CB5CDDEBF7DBB2DAAA159";
    attribute INIT_07 of inst : label is "CEA4884CFB9FFEC7EF249CC9295ABABB11454513E1FFACF8FFEB3E3FFAD5377A";
    attribute INIT_08 of inst : label is "D9359A4A3408EC65914BB0A13C644BF6E44CCBFC003C002C52EDFB72266446C8";
    attribute INIT_09 of inst : label is "08BAABAB47625ECECC962D5078B55C38720204A3F7220A1B334088464496D345";
    attribute INIT_0A of inst : label is "AEBAE1534C298532A645142D5716ABEB14907F483FA41FD20FEBB19554CA2C25";
    attribute INIT_0B of inst : label is "5819141A6450699141A6450710B40CA74E9C1E9D3A707F5A74E9D1E9D3A747F5";
    attribute INIT_0C of inst : label is "948D390EEB0090C2C090CC2CAD4AA4561740B5C4EE4AEB2EC0F13B3FF2C44466";
    attribute INIT_0D of inst : label is "7755B8EC930D86C6D22110812626270B06E3B23BBBB8DC765BEEEEE2B71D8538";
    attribute INIT_0E of inst : label is "EAA1820044009CFD8AFFFFFF0004FFFFFFF00000000FFF00F5AB76AD00B71D92";
    attribute INIT_0F of inst : label is "0F389ADD755038909853572D80584092A9CA644452D62F5555AB6592AFF53E59";
    attribute INIT_10 of inst : label is "BA240D1A25E7AF30DDDDFF83DF32F7FDFBFEFFDFF9F7AD6F0DF5ADEB0DB5ADEF";
    attribute INIT_11 of inst : label is "C2D88385C0023BE2C2438B24B1A91A894C36B62423421B94891304111737C91A";
    attribute INIT_12 of inst : label is "6D1957831162A5188E5B32990C452224818006085E486002986C56114000070A";
    attribute INIT_13 of inst : label is "2DC185B83F465B6BB0F0FBAD54CB868D2C813C370000000034C132689948D024";
    attribute INIT_14 of inst : label is "E687271049000BA9008AA1D2B0A252884A2147000521002120DB830B72616E4C";
    attribute INIT_15 of inst : label is "6AC34994340C5D0721068994A4C2401A34E1400000000636415BC512E9D142EB";
    attribute INIT_16 of inst : label is "F800487A208002989A00000D124C4DA952DA1B52B62FB25295524C24524982D8";
    attribute INIT_17 of inst : label is "9EE73DCF73DCF73CE639CE7398C7318E63AC068E80907B4CCBB2444D2483FF87";
    attribute INIT_18 of inst : label is "D5C81D00000000000000000000000040400050800510A00344C80344C2022F13";
    attribute INIT_19 of inst : label is "8BDA14C5ED0A602AA9AAC772B340975CB8EE3971EDBD6F50B4E07121A9404CD2";
    attribute INIT_1A of inst : label is "8351A31A4404CD34000000011F1F1F6363EB1EF0B7A3CBEFFFD199C320D6BC2D";
    attribute INIT_1B of inst : label is "280000220010DA85D31694946B1A25090246CDB11DA782994CA6532982A86A1A";
    attribute INIT_1C of inst : label is "2AA3AA7382A8EA9C50AA8EA9D340AA66DB3C17ED92E6F65B4E4EE596369824C6";
    attribute INIT_1D of inst : label is "400004104104115140000410410418E09003F88EA9DC271DD2271CE0AA3AA714";
    attribute INIT_1E of inst : label is "0000000020202020000000004A40A82A084A288A088045055514155450555151";
    attribute INIT_1F of inst : label is "A00C030A86B058818B30B3564C0E0DD7044440A1455155554515111222222222";
    attribute INIT_20 of inst : label is "899F8F6B75BB4945A48001290044B122119813A324BBFEFEE5008421284A1084";
    attribute INIT_21 of inst : label is "4000A048192902D40C8140C96AF219025D40C011CE4899F5F6AF018025FA0640";
    attribute INIT_22 of inst : label is "000002A2035C2493B812481626524892641524C82924E880D2429092E630ABC2";
    attribute INIT_23 of inst : label is "FF740FFFFFBFFFFDF0000400AA02AA02AB0005035555540000000035444D0000";
    attribute INIT_24 of inst : label is "873CDE79471479ECF38404FB6DA7DE0E7FEFFF9E0FFFFEFFFD07DFEEFFFFC3EF";
    attribute INIT_25 of inst : label is "3829EEBAD522BAFF02BBEB0F7D75F4DF36FBCD7CB8C3FFF7EEFF5F5FDBFBDFF0";
    attribute INIT_26 of inst : label is "079C0FF9FEBBFFF400CB7EFFC3F8FF8B7FBF8FF77FB9E0F3CE0051E78C00A0CF";
    attribute INIT_27 of inst : label is "7FFFFFFFF13F07F13F07F13F07F0FFF7FFBFF7FFBFF7FFF83FFDF03C03A00210";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "2CBB2BF35FA1FFFF6B4D83E4AC8696D07666FA7FFFFFFFFFF8FFE82155016D8B";
    attribute INIT_01 of inst : label is "04B44CCB4A54A964A44924926492E1009AA82B5AE95B55AAFFFFFFF86BF92DDD";
    attribute INIT_02 of inst : label is "1AD6D10D3036C30D30364528A516A29452A014EDD5DBF6A74AE52B6969008401";
    attribute INIT_03 of inst : label is "50AAEBCE900000490209918209204132B4412408264608248104CAC15ADB0076";
    attribute INIT_04 of inst : label is "E132C2A929961D48822D3A652B3657AABA65855202F3A6709CA9AB4E9B4B4555";
    attribute INIT_05 of inst : label is "77222C821108442110825214A527C8C821AA915544DC4069EAA6CB28132C3A94";
    attribute INIT_06 of inst : label is "4924E6AF2CE92D5C88B22A9AB24925357967496EE4459154D5924929ABCB3A4B";
    attribute INIT_07 of inst : label is "CA948A554B9908E642A4DCCB2958A8AB104541113739644D4E59135396475356";
    attribute INIT_08 of inst : label is "CB2C9E492508A3249949908165654992264CE8E6A826A8265264C9132654624C";
    attribute INIT_09 of inst : label is "0C88A889351A4A0ECCD6A8208895474E9240008273524E88D25088565493D154";
    attribute INIT_0A of inst : label is "49249B3289112224448C60255112A8D2689299494CA4A652532B719AA8CDA832";
    attribute INIT_0B of inst : label is "523B1458EC5163B1458EC51638A03244891231122458D9144891231122458D91";
    attribute INIT_0C of inst : label is "AC2BE84EEB802006C020106C260A3112B2408584ED484E04E09B28A49AD55555";
    attribute INIT_0D of inst : label is "DB55A2F3938DC6E6D02010010606061B068BCE313B8BD179C4C4EE2EA45E6BEA";
    attribute INIT_0E of inst : label is "2AA0135566AACE701FFF00000000FF000FFFFF96000FFFFF055A956814D45E72";
    attribute INIT_0F of inst : label is "A5019294BAA0D9211021436510DA4992AC546555528830FF3DFB5506420240A3";
    attribute INIT_10 of inst : label is "0A0806014086843807C52983653294E7289392524CE529CAA4E7294EA4A7294A";
    attribute INIT_11 of inst : label is "03822D86C0403B329243AB2630400C194E373608418017CC8608042994366104";
    attribute INIT_12 of inst : label is "2641463B5A748508885733198445BBAC820808201F0080010002080080021001";
    attribute INIT_13 of inst : label is "0451808A3006DBABB2C0804C45DB141AEA3030080000000000093A6820D82008";
    attribute INIT_14 of inst : label is "C4024390008388B82B14CDD529AAD6AB5AFD61A00A0228280008B3011460228C";
    attribute INIT_15 of inst : label is "30009B20086C6E24C126820DA0E082041109500000000000B84C16A223A26279";
    attribute INIT_16 of inst : label is "FFFFB079556A8004209FFC1000000040E7002081C02C90469F52DA4E7E5B4A4C";
    attribute INIT_17 of inst : label is "484290A5294A5294A521485294A5290A52A40329006724CAD990054B6003FC7F";
    attribute INIT_18 of inst : label is "56D0220000000000000000FFFFFF7F041FBFA41FDA40402F8810178804000009";
    attribute INIT_19 of inst : label is "51CE0120E701902A88A883209201264F90641B20E7294E700B61B24146001244";
    attribute INIT_1A of inst : label is "02A5040D200124C6000000008E8E8A6E514E8E5018C1A929CE7010602A439402";
    attribute INIT_1B of inst : label is "13FFFF956A804C95B60728149A04180601826F045D9604924924924905405014";
    attribute INIT_1C of inst : label is "AAA0A82380A82A0802AA82A09283245492A805C924AE84D2EA94AD3476B4CDCD";
    attribute INIT_1D of inst : label is "444510441041011044451044104108A00AA8A082A09A2208822208E02A0A8200";
    attribute INIT_1E of inst : label is "202020202020202020202020406004010008AA8A088055055554155550555110";
    attribute INIT_1F of inst : label is "40520972C1D86D31177F0062288269A204504201111511115555555202020202";
    attribute INIT_20 of inst : label is "A99279681FBB8B4D84C92843184CB9841391369B64CA739E888981C0501C0701";
    attribute INIT_21 of inst : label is "E2A8EC7B1B2B82DD8DC1D8D96E371B8267D8DC150D4A992696E371B8252EC6E0";
    attribute INIT_22 of inst : label is "0000028627C56D860E3EDE74AD74DA94EE3F69DC7564A189F4C2B85329BCA8C2";
    attribute INIT_23 of inst : label is "2275D000AAEAAA0200000C0132033203320030602AAA2AAA8AAAA04200000000";
    attribute INIT_24 of inst : label is "000000008208000000001A80924C21F6002000000480000000F8000100148210";
    attribute INIT_25 of inst : label is "003E114F9555453FFD443C028AAA0B20C9063A83060000000000202000002000";
    attribute INIT_26 of inst : label is "F8020006596402F7DE36DB00000704708004700CA4580000020000C094000380";
    attribute INIT_27 of inst : label is "7FFFFFFFE03F07F03F07F03F07F0000800400800400801040081F7C3FC534D27";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "248921294484FFFFE13F98120210721989123FFFFFFFFFFFF9FFF80011408A38";
    attribute INIT_01 of inst : label is "FB0672306387301837B6DB6D9B6D0C92618D942105C87083FFFFFFF92894244C";
    attribute INIT_02 of inst : label is "E3296616400974164009ECE59CB39672CE56C712062408587318E085849277BC";
    attribute INIT_03 of inst : label is "1288C470E0000395B50E623C70B6A1CCC38E16D4399871C2DA87331EC9046CC8";
    attribute INIT_04 of inst : label is "80CD1D2E0668E976C8E5A99884C18822319A3A5C013C38C0674E06F4EA748111";
    attribute INIT_05 of inst : label is "31CDD34BEE2FB8BEE6491CC731D83735D855FAAAEAF37626555934CC0CD1C2E7";
    attribute INIT_06 of inst : label is "B6DB5A03DF0EDCC7374DC0E08DB6D8D01EF876E639BA6E07046DB6C680F7C3B7";
    attribute INIT_07 of inst : label is "30C77784F46671199C3B2734D6A02828DBAC6EBEC3C61BB07186EC3C61BA1C11";
    attribute INIT_08 of inst : label is "34C365ADB1F730DB662E62041A9AB6EDD9734F1955D955D98B9B76ECB9A79DB3";
    attribute INIT_09 of inst : label is "32F70F75A183337133282DD8772AB870EB7BDE7D801D74EC1B1F7129AB6C1E27";
    attribute INIT_0A of inst : label is "2CB2C48C44C89913227093CAAEE5574B90D8E66C7336399B1CD496655B322CCD";
    attribute INIT_0B of inst : label is "5BC4061F10187C4061F10187C734CB224489C089122706E224489C089122706E";
    attribute INIT_0C of inst : label is "8C9921392479500139502813DA61C0EC3D82DA1310B332334360CD1B65044444";
    attribute INIT_0D of inst : label is "DAABA0F4FC3219093B81C0C4B83838041E83D3E88880D07A72A22203341E9920";
    attribute INIT_0E of inst : label is "15670CAAD955B5B140F0FFFFFFFF00FFFFFF6969FFF000000DAB56AD2A341E9E";
    attribute INIT_0F of inst : label is "39846C63355098F3D8DE0C1B4E2595E55EB398445AF6C95515AB0593A2104183";
    attribute INIT_10 of inst : label is "2044150DD63831C438B8C68C18CC631AD76C6D8DB358C6B43B5AC6343B18C630";
    attribute INIT_11 of inst : label is "FDEC1984C984C4CC5D9C0CD8E2A02A0670C8485404431023110D92C661C90E22";
    attribute INIT_12 of inst : label is "31661843238758277589CD6613BA22233DF6F7DFC0FF7DFEFF7DF7DF77FDEFBE";
    attribute INIT_13 of inst : label is "800E1001C098A40C4CD2D8B000042E792C9DC054000000005965C38150215054";
    attribute INIT_14 of inst : label is "96CC3CC7DF78335EC94D3BCEB602C81F202CB00F858D8787A9001C2003840070";
    attribute INIT_15 of inst : label is "88244410444C4D36A1B815023705412A1A941800000002035ABA41D00C1D3F96";
    attribute INIT_16 of inst : label is "0000007AAA955FFBDF4001EFDFEFEFBF18FBDF7E3F80CB0840182191010439B0";
    attribute INIT_17 of inst : label is "695AD2B5AD6B5AD6B5AD695AD6B5AD6B5ADA428AC811C220266B10608FFFFC78";
    attribute INIT_18 of inst : label is "8CDCF1000000000000000000000000FBE0005BE005BFBFC077EFE077FBFBFFED";
    attribute INIT_19 of inst : label is "26B0429B58204C9575571CC70B4AB9B06398E0C718C63182066131E5F1040B6B";
    attribute INIT_1A of inst : label is "C3579270B042B63800000000747471838E307182170E16C631820384038C6085";
    attribute INIT_1B of inst : label is "E800002A955962C608591EC3C30A5415054343D8224682592C964B2582AC6B1A";
    attribute INIT_1C of inst : label is "2AAAAAA280AAAAA880AAAAAA9B1EDB66DB39B70DB6C6C61B4ED8C1C7D363A340";
    attribute INIT_1D of inst : label is "404100441041015140410044104109A02002AA8AAA88A22882A228A02AAAAA20";
    attribute INIT_1E of inst : label is "A8A8A8A8A8A8A8A8A8A8A8A8C4405415042AAA8A085500500001400005000151";
    attribute INIT_1F of inst : label is "240B05AB4068964321D9213BF20B928C0455400155151515551515162AAAAAAA";
    attribute INIT_20 of inst : label is "0E6C8EC4E1E6B0633306779CEF6366325EB28CC6DB318C62245710A429024090";
    attribute INIT_21 of inst : label is "51571785E0D91D82F48E2F06C1D2E84D982F42613070E6C9EC1D0E84D8D17A07";
    attribute INIT_22 of inst : label is "000009DD5D08CB5871E12316384B20EB99E4D733C1D2F7574B2D919DBD16E75C";
    attribute INIT_23 of inst : label is "0076200000400002100006003C003C003DC1CF9F55555555555557BDF7FFF000";
    attribute INIT_24 of inst : label is "0C01200082080201000C1280105000018014181200007D0002F820117C100250";
    attribute INIT_25 of inst : label is "000200001588103F000041082010470820000000430008081100A8A024042000";
    attribute INIT_26 of inst : label is "00800076820800F42B208360008820F68F60800892500001C000200310004380";
    attribute INIT_27 of inst : label is "7FFFFFFC00000000000000000000106B8C78CB0C7CCB09240001F803000CB0C8";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "201801110400FFFFC03F90000402205900007FFFFFFFFFFFF9FFF80011000831";
    attribute INIT_01 of inst : label is "A012044122041A2116000000200025B6C30DB8002C812001FFFFFFF820880040";
    attribute INIT_02 of inst : label is "C231C01C0011C01C00118841082104208436C200440000604120410D0DB6D294";
    attribute INIT_03 of inst : label is "1288844080000220A50802104414A100C208C294201841105284011880082DD0";
    attribute INIT_04 of inst : label is "8080112884008946484488018C0218222100205101B12240644886C48A448111";
    attribute INIT_05 of inst : label is "3110044900240090024B104431024005115572AA8A9070141550000408011282";
    attribute INIT_06 of inst : label is "000000070C0808C4401110809000020038604046220088040480000001C30202";
    attribute INIT_07 of inst : label is "00C4420C404040101020440118A030314A082828130022044008813002201012";
    attribute INIT_08 of inst : label is "0104042590801500082802042080800003400C01550155020A000001A0063004";
    attribute INIT_09 of inst : label is "0640040480A9616200682511402AA04089294A50001140E54908010808010804";
    attribute INIT_0A of inst : label is "24924810444889112220160AA805544918488024401220091014A00558022411";
    attribute INIT_0B of inst : label is "4988061620185880616201858C140B2244888089122208022448880891222080";
    attribute INIT_0C of inst : label is "8819003A00B9500239502823026311802006CC3600C30630000904000D044444";
    attribute INIT_0D of inst : label is "D8ABA0B2F82010103B0180C0B03030081A82CBC88880D0597222220394165900";
    attribute INIT_0E of inst : label is "154400AA815500100AF0FFFFFFFFFF0000000000000000F008A142850A34165C";
    attribute INIT_0F of inst : label is "208C800B255090F3C81800235C4615055DB200444A46195514A9048222024182";
    attribute INIT_10 of inst : label is "0044150DD630318C626000004280000204000000044000042042008420000000";
    attribute INIT_11 of inst : label is "0700390489C580105E080802E22022082080404404431044110DB6D081802E22";
    attribute INIT_12 of inst : label is "117018F232244020040901009002222400000000000000000000000000000000";
    attribute INIT_13 of inst : label is "8004100080B080880C9250A000880A79041D8054000000004B6C890150415054";
    attribute INIT_14 of inst : label is "A2803080000000700B0C390E9C02801E0028E000000000000900082001040020";
    attribute INIT_15 of inst : label is "A825485044484912A0B015041625432A08B818000000026C72770EC57A9EC410";
    attribute INIT_16 of inst : label is "FFFFB7800000000000000000000000000000000001044B000010408202081004";
    attribute INIT_17 of inst : label is "2B5A5694A5294A5294A5295A52B4A5694AE24088C8510A40400B00410007FC7F";
    attribute INIT_18 of inst : label is "0C9CF5000000000000000000000000000000000000000000000000000000002D";
    attribute INIT_19 of inst : label is "700040B800205C85415410046142A0008200810400100402064121E4F5040B22";
    attribute INIT_1A of inst : label is "C1528245B042B2A200000000C4C0C0021800C002044838000422022402200081";
    attribute INIT_1B of inst : label is "88000000000B22C410D91EC3C90A541505410600406482492492492482AC2B0A";
    attribute INIT_1C of inst : label is "A220200A2A8808022A88808039B8E33249139344924642490448449301822444";
    attribute INIT_1D of inst : label is "1514551145145404151455114514588A8AA88020802A0882AA08828AA202008A";
    attribute INIT_1E of inst : label is "0202020202020202020202024055014050080828A85555555555555555555404";
    attribute INIT_1F of inst : label is "240B0CABC0781C0132092139E009028E05004001015151510151515200000000";
    attribute INIT_20 of inst : label is "080098058D808124304656B4AD2408A230B31040004001000054102409024090";
    attribute INIT_21 of inst : label is "0154362D81000006C0006C0803000100226C0801004080098030201000136040";
    attribute INIT_22 of inst : label is "000009905100085CC58B21122059208A018D140311126414593000119C124400";
    attribute INIT_23 of inst : label is "3F8BF0000000000210000801C003C003C0000000000000000000000000000000";
    attribute INIT_24 of inst : label is "000000000200000000001280104000000004181200007C0000F800007C100210";
    attribute INIT_25 of inst : label is "0002000AEA8C0AC0AC0041000010470820000000000000000000082000000000";
    attribute INIT_26 of inst : label is "0000003682083F0BF8208360000820F20F208008925000018208200304104380";
    attribute INIT_27 of inst : label is "7FFFFFFC0000000000000000000010430C38C30C3CC3092400FE0FC300000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
