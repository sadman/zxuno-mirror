-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e3",
     9 => x"c4080b0b",
    10 => x"80e3c808",
    11 => x"0b0b80e3",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e3cc0c0b",
    16 => x"0b80e3c8",
    17 => x"0c0b0b80",
    18 => x"e3c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80ddf0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e3c470",
    57 => x"80edfc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51b18c",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e3",
    65 => x"d40c9f0b",
    66 => x"80e3d80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e3d808ff",
    70 => x"0580e3d8",
    71 => x"0c80e3d8",
    72 => x"088025e8",
    73 => x"3880e3d4",
    74 => x"08ff0580",
    75 => x"e3d40c80",
    76 => x"e3d40880",
    77 => x"25d03880",
    78 => x"0b80e3d8",
    79 => x"0c800b80",
    80 => x"e3d40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e3d408",
   100 => x"25913882",
   101 => x"c82d80e3",
   102 => x"d408ff05",
   103 => x"80e3d40c",
   104 => x"838a0480",
   105 => x"e3d40880",
   106 => x"e3d80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e3d408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e3d80881",
   116 => x"0580e3d8",
   117 => x"0c80e3d8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e3d8",
   121 => x"0c80e3d4",
   122 => x"08810580",
   123 => x"e3d40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e3",
   128 => x"d8088105",
   129 => x"80e3d80c",
   130 => x"80e3d808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e3d8",
   134 => x"0c80e3d4",
   135 => x"08810580",
   136 => x"e3d40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e3dc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e3dc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e3",
   177 => x"dc088407",
   178 => x"80e3dc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80e0",
   183 => x"b00c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e3dc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e3",
   208 => x"c40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"a00bec0c",
  1093 => x"86c72d86",
  1094 => x"c72d86c7",
  1095 => x"2d86c72d",
  1096 => x"86c72d86",
  1097 => x"c72d86c7",
  1098 => x"2d86c72d",
  1099 => x"86c72d86",
  1100 => x"c72d86c7",
  1101 => x"2d86c72d",
  1102 => x"86c72d86",
  1103 => x"c72d86c7",
  1104 => x"2d86c72d",
  1105 => x"86c72d86",
  1106 => x"c72d86c7",
  1107 => x"2d86c72d",
  1108 => x"86c72d86",
  1109 => x"c72d86c7",
  1110 => x"2d86c72d",
  1111 => x"86c72d86",
  1112 => x"c72d86c7",
  1113 => x"2d86c72d",
  1114 => x"86c72d86",
  1115 => x"c72d86c7",
  1116 => x"2d86c72d",
  1117 => x"86c72d86",
  1118 => x"c72d86c7",
  1119 => x"2d86c72d",
  1120 => x"86c72d86",
  1121 => x"c72d86c7",
  1122 => x"2d86c72d",
  1123 => x"86c72d86",
  1124 => x"c72d86c7",
  1125 => x"2d86c72d",
  1126 => x"86c72d86",
  1127 => x"c72d86c7",
  1128 => x"2d86c72d",
  1129 => x"86c72d86",
  1130 => x"c72d86c7",
  1131 => x"2d86c72d",
  1132 => x"86c72d86",
  1133 => x"c72d86c7",
  1134 => x"2d86c72d",
  1135 => x"86c72d86",
  1136 => x"c72d86c7",
  1137 => x"2d86c72d",
  1138 => x"86c72d86",
  1139 => x"c72d86c7",
  1140 => x"2d86c72d",
  1141 => x"86c72d86",
  1142 => x"c72d86c7",
  1143 => x"2d86c72d",
  1144 => x"86c72d86",
  1145 => x"c72d86c7",
  1146 => x"2d86c72d",
  1147 => x"86c72d86",
  1148 => x"c72d86c7",
  1149 => x"2d86c72d",
  1150 => x"86c72d86",
  1151 => x"c72d86c7",
  1152 => x"2d86c72d",
  1153 => x"86c72d86",
  1154 => x"c72d86c7",
  1155 => x"2d86c72d",
  1156 => x"86c72d86",
  1157 => x"c72d86c7",
  1158 => x"2d86c72d",
  1159 => x"86c72d86",
  1160 => x"c72d86c7",
  1161 => x"2d86c72d",
  1162 => x"86c72d86",
  1163 => x"c72d86c7",
  1164 => x"2d86c72d",
  1165 => x"86c72d86",
  1166 => x"c72d86c7",
  1167 => x"2d86c72d",
  1168 => x"86c72d86",
  1169 => x"c72d86c7",
  1170 => x"2d86c72d",
  1171 => x"86c72d86",
  1172 => x"c72d86c7",
  1173 => x"2d86c72d",
  1174 => x"86c72d86",
  1175 => x"c72d86c7",
  1176 => x"2d86c72d",
  1177 => x"86c72d86",
  1178 => x"c72d86c7",
  1179 => x"2d86c72d",
  1180 => x"86c72d86",
  1181 => x"c72d86c7",
  1182 => x"2d86c72d",
  1183 => x"86c72d86",
  1184 => x"c72d86c7",
  1185 => x"2d86c72d",
  1186 => x"86c72d86",
  1187 => x"c72d86c7",
  1188 => x"2d86c72d",
  1189 => x"86c72d86",
  1190 => x"c72d86c7",
  1191 => x"2d86c72d",
  1192 => x"86c72d86",
  1193 => x"c72d86c7",
  1194 => x"2d86c72d",
  1195 => x"86c72d86",
  1196 => x"c72d86c7",
  1197 => x"2d86c72d",
  1198 => x"86c72d86",
  1199 => x"c72d86c7",
  1200 => x"2d86c72d",
  1201 => x"86c72d86",
  1202 => x"c72d86c7",
  1203 => x"2d86c72d",
  1204 => x"86c72d86",
  1205 => x"c72d86c7",
  1206 => x"2d86c72d",
  1207 => x"86c72d86",
  1208 => x"c72d86c7",
  1209 => x"2d86c72d",
  1210 => x"86c72d86",
  1211 => x"c72d86c7",
  1212 => x"2d86c72d",
  1213 => x"86c72d86",
  1214 => x"c72d86c7",
  1215 => x"2d86c72d",
  1216 => x"86c72d86",
  1217 => x"c72d86c7",
  1218 => x"2d86c72d",
  1219 => x"86c72d86",
  1220 => x"c72d86c7",
  1221 => x"2d86c72d",
  1222 => x"86c72d86",
  1223 => x"c72d86c7",
  1224 => x"2d86c72d",
  1225 => x"86c72d86",
  1226 => x"c72d86c7",
  1227 => x"2d86c72d",
  1228 => x"86c72d86",
  1229 => x"c72d86c7",
  1230 => x"2d86c72d",
  1231 => x"86c72d86",
  1232 => x"c72d86c7",
  1233 => x"2d86c72d",
  1234 => x"86c72d86",
  1235 => x"c72d86c7",
  1236 => x"2d86c72d",
  1237 => x"86c72d86",
  1238 => x"c72d86c7",
  1239 => x"2d86c72d",
  1240 => x"86c72d86",
  1241 => x"c72d86c7",
  1242 => x"2d86c72d",
  1243 => x"86c72d86",
  1244 => x"c72d86c7",
  1245 => x"2d86c72d",
  1246 => x"86c72d86",
  1247 => x"c72d86c7",
  1248 => x"2d86c72d",
  1249 => x"86c72d86",
  1250 => x"c72d86c7",
  1251 => x"2d86c72d",
  1252 => x"86c72d86",
  1253 => x"c72d86c7",
  1254 => x"2d86c72d",
  1255 => x"86c72d86",
  1256 => x"c72d86c7",
  1257 => x"2d86c72d",
  1258 => x"86c72d86",
  1259 => x"c72d86c7",
  1260 => x"2d86c72d",
  1261 => x"86c72d86",
  1262 => x"c72d86c7",
  1263 => x"2d86c72d",
  1264 => x"86c72d86",
  1265 => x"c72d86c7",
  1266 => x"2d86c72d",
  1267 => x"86c72d86",
  1268 => x"c72d86c7",
  1269 => x"2d86c72d",
  1270 => x"86c72d86",
  1271 => x"c72d86c7",
  1272 => x"2d86c72d",
  1273 => x"86c72d86",
  1274 => x"c72d86c7",
  1275 => x"2d86c72d",
  1276 => x"86c72d86",
  1277 => x"c72d86c7",
  1278 => x"2d86c72d",
  1279 => x"86c72d86",
  1280 => x"c72d86c7",
  1281 => x"2d86c72d",
  1282 => x"86c72d86",
  1283 => x"c72d86c7",
  1284 => x"2d86c72d",
  1285 => x"86c72d86",
  1286 => x"c72d86c7",
  1287 => x"2d86c72d",
  1288 => x"86c72d86",
  1289 => x"c72d86c7",
  1290 => x"2d86c72d",
  1291 => x"86c72d86",
  1292 => x"c72d86c7",
  1293 => x"2d86c72d",
  1294 => x"86c72d86",
  1295 => x"c72d86c7",
  1296 => x"2d86c72d",
  1297 => x"86c72d86",
  1298 => x"c72d86c7",
  1299 => x"2d86c72d",
  1300 => x"86c72d86",
  1301 => x"c72d86c7",
  1302 => x"2d86c72d",
  1303 => x"86c72d86",
  1304 => x"c72d86c7",
  1305 => x"2d86c72d",
  1306 => x"86c72d86",
  1307 => x"c72d86c7",
  1308 => x"2d86c72d",
  1309 => x"86c72d86",
  1310 => x"c72d86c7",
  1311 => x"2d86c72d",
  1312 => x"86c72d86",
  1313 => x"c72d86c7",
  1314 => x"2d86c72d",
  1315 => x"86c72d86",
  1316 => x"c72d86c7",
  1317 => x"2d86c72d",
  1318 => x"86c72d86",
  1319 => x"c72d86c7",
  1320 => x"2d86c72d",
  1321 => x"86c72d86",
  1322 => x"c72d86c7",
  1323 => x"2d86c72d",
  1324 => x"86c72d86",
  1325 => x"c72d86c7",
  1326 => x"2d86c72d",
  1327 => x"86c72d86",
  1328 => x"c72d86c7",
  1329 => x"2d86c72d",
  1330 => x"86c72d86",
  1331 => x"c72d86c7",
  1332 => x"2d86c72d",
  1333 => x"86c72d86",
  1334 => x"c72d86c7",
  1335 => x"2d86c72d",
  1336 => x"86c72d86",
  1337 => x"c72d86c7",
  1338 => x"2d86c72d",
  1339 => x"86c72d86",
  1340 => x"c72d86c7",
  1341 => x"2d86c72d",
  1342 => x"86c72d86",
  1343 => x"c72d86c7",
  1344 => x"2d86c72d",
  1345 => x"86c72d86",
  1346 => x"c72d86c7",
  1347 => x"2d86c72d",
  1348 => x"86c72d86",
  1349 => x"c72d86c7",
  1350 => x"2d86c72d",
  1351 => x"86c72d86",
  1352 => x"c72d86c7",
  1353 => x"2d86c72d",
  1354 => x"86c72d86",
  1355 => x"c72d86c7",
  1356 => x"2d86c72d",
  1357 => x"86c72d86",
  1358 => x"c72d86c7",
  1359 => x"2d86c72d",
  1360 => x"86c72d86",
  1361 => x"c72d86c7",
  1362 => x"2d86c72d",
  1363 => x"86c72d86",
  1364 => x"c72d86c7",
  1365 => x"2d86c72d",
  1366 => x"86c72d86",
  1367 => x"c72d86c7",
  1368 => x"2d86c72d",
  1369 => x"86c72d86",
  1370 => x"c72d86c7",
  1371 => x"2d86c72d",
  1372 => x"86c72d86",
  1373 => x"c72d86c7",
  1374 => x"2d86c72d",
  1375 => x"86c72d86",
  1376 => x"c72d86c7",
  1377 => x"2d86c72d",
  1378 => x"86c72d86",
  1379 => x"c72d86c7",
  1380 => x"2d86c72d",
  1381 => x"86c72d86",
  1382 => x"c72d86c7",
  1383 => x"2d86c72d",
  1384 => x"86c72d86",
  1385 => x"c72d86c7",
  1386 => x"2d86c72d",
  1387 => x"86c72d86",
  1388 => x"c72d86c7",
  1389 => x"2d86c72d",
  1390 => x"86c72d86",
  1391 => x"c72d86c7",
  1392 => x"2d86c72d",
  1393 => x"86c72d86",
  1394 => x"c72d86c7",
  1395 => x"2d86c72d",
  1396 => x"86c72d86",
  1397 => x"c72d86c7",
  1398 => x"2d86c72d",
  1399 => x"86c72d86",
  1400 => x"c72d86c7",
  1401 => x"2d86c72d",
  1402 => x"86c72d86",
  1403 => x"c72d86c7",
  1404 => x"2d86c72d",
  1405 => x"86c72d86",
  1406 => x"c72d86c7",
  1407 => x"2d86c72d",
  1408 => x"86c72d86",
  1409 => x"c72d86c7",
  1410 => x"2d86c72d",
  1411 => x"86c72d86",
  1412 => x"c72d86c7",
  1413 => x"2d86c72d",
  1414 => x"86c72d86",
  1415 => x"c72d86c7",
  1416 => x"2d86c72d",
  1417 => x"86c72d86",
  1418 => x"c72d86c7",
  1419 => x"2d86c72d",
  1420 => x"86c72d86",
  1421 => x"c72d86c7",
  1422 => x"2d86c72d",
  1423 => x"86c72d86",
  1424 => x"c72d86c7",
  1425 => x"2d86c72d",
  1426 => x"86c72d86",
  1427 => x"c72d86c7",
  1428 => x"2d86c72d",
  1429 => x"86c72d86",
  1430 => x"c72d86c7",
  1431 => x"2d86c72d",
  1432 => x"86c72d86",
  1433 => x"c72d86c7",
  1434 => x"2d86c72d",
  1435 => x"86c72d86",
  1436 => x"c72d86c7",
  1437 => x"2d86c72d",
  1438 => x"86c72d86",
  1439 => x"c72d86c7",
  1440 => x"2d86c72d",
  1441 => x"86c72d86",
  1442 => x"c72d86c7",
  1443 => x"2d86c72d",
  1444 => x"86c72d86",
  1445 => x"c72d86c7",
  1446 => x"2d86c72d",
  1447 => x"86c72d86",
  1448 => x"c72d86c7",
  1449 => x"2d86c72d",
  1450 => x"86c72d86",
  1451 => x"c72d86c7",
  1452 => x"2d86c72d",
  1453 => x"86c72d86",
  1454 => x"c72d86c7",
  1455 => x"2d86c72d",
  1456 => x"86c72d86",
  1457 => x"c72d86c7",
  1458 => x"2d86c72d",
  1459 => x"86c72d86",
  1460 => x"c72d86c7",
  1461 => x"2d86c72d",
  1462 => x"86c72d86",
  1463 => x"c72d86c7",
  1464 => x"2d86c72d",
  1465 => x"86c72d86",
  1466 => x"c72d86c7",
  1467 => x"2d86c72d",
  1468 => x"86c72d86",
  1469 => x"c72d86c7",
  1470 => x"2d86c72d",
  1471 => x"86c72d86",
  1472 => x"c72d86c7",
  1473 => x"2d86c72d",
  1474 => x"86c72d86",
  1475 => x"c72d86c7",
  1476 => x"2d86c72d",
  1477 => x"86c72d86",
  1478 => x"c72d86c7",
  1479 => x"2d86c72d",
  1480 => x"86c72d86",
  1481 => x"c72d86c7",
  1482 => x"2d86c72d",
  1483 => x"86c72d86",
  1484 => x"c72d86c7",
  1485 => x"2d86c72d",
  1486 => x"86c72d86",
  1487 => x"c72d86c7",
  1488 => x"2d86c72d",
  1489 => x"86c72d86",
  1490 => x"c72d86c7",
  1491 => x"2d86c72d",
  1492 => x"86c72d86",
  1493 => x"c72d86c7",
  1494 => x"2d86c72d",
  1495 => x"86c72d86",
  1496 => x"c72d86c7",
  1497 => x"2d86c72d",
  1498 => x"86c72d86",
  1499 => x"c72d86c7",
  1500 => x"2d86c72d",
  1501 => x"86c72d86",
  1502 => x"c72d86c7",
  1503 => x"2d86c72d",
  1504 => x"86c72d86",
  1505 => x"c72d86c7",
  1506 => x"2d86c72d",
  1507 => x"86c72d86",
  1508 => x"c72d86c7",
  1509 => x"2d86c72d",
  1510 => x"86c72d86",
  1511 => x"c72d86c7",
  1512 => x"2d86c72d",
  1513 => x"86c72d86",
  1514 => x"c72d86c7",
  1515 => x"2d86c72d",
  1516 => x"86c72d86",
  1517 => x"c72d86c7",
  1518 => x"2d86c72d",
  1519 => x"86c72d86",
  1520 => x"c72d86c7",
  1521 => x"2d86c72d",
  1522 => x"86c72d86",
  1523 => x"c72d86c7",
  1524 => x"2d86c72d",
  1525 => x"0402dc05",
  1526 => x"0d8059a2",
  1527 => x"902d810b",
  1528 => x"ec0c7a52",
  1529 => x"80e3e051",
  1530 => x"80d4bd2d",
  1531 => x"80e3c408",
  1532 => x"792e80f7",
  1533 => x"3880e3e4",
  1534 => x"0870f80c",
  1535 => x"79ff1256",
  1536 => x"59557379",
  1537 => x"2e8b3881",
  1538 => x"1874812a",
  1539 => x"555873f7",
  1540 => x"38f71858",
  1541 => x"81598075",
  1542 => x"2580d038",
  1543 => x"77527351",
  1544 => x"84a82d80",
  1545 => x"e4b45280",
  1546 => x"e3e05180",
  1547 => x"d7932d80",
  1548 => x"e3c40880",
  1549 => x"2e9b3880",
  1550 => x"e4b45783",
  1551 => x"fc567670",
  1552 => x"84055808",
  1553 => x"e80cfc16",
  1554 => x"56758025",
  1555 => x"f138b0d9",
  1556 => x"0480e3c4",
  1557 => x"08598480",
  1558 => x"5580e3e0",
  1559 => x"5180d6e2",
  1560 => x"2dfc8015",
  1561 => x"81155555",
  1562 => x"b0960484",
  1563 => x"0bec0c78",
  1564 => x"802e8838",
  1565 => x"80e0b451",
  1566 => x"b0ff0480",
  1567 => x"e19451b8",
  1568 => x"c12d7880",
  1569 => x"e3c40c02",
  1570 => x"a4050d04",
  1571 => x"02f0050d",
  1572 => x"840bec0c",
  1573 => x"b5fe2db2",
  1574 => x"b32d81f9",
  1575 => x"2d8352b5",
  1576 => x"e12d8151",
  1577 => x"858d2dff",
  1578 => x"12527180",
  1579 => x"25f13884",
  1580 => x"0bec0c80",
  1581 => x"dee45186",
  1582 => x"a02d80ca",
  1583 => x"dd2d80e3",
  1584 => x"c408802e",
  1585 => x"80d638af",
  1586 => x"d55180dd",
  1587 => x"ea2d80e0",
  1588 => x"b451b8c1",
  1589 => x"2db6a02d",
  1590 => x"b2bf2db8",
  1591 => x"d42d80e0",
  1592 => x"c80b80f5",
  1593 => x"2d80e280",
  1594 => x"08708106",
  1595 => x"54555371",
  1596 => x"802e8538",
  1597 => x"72810753",
  1598 => x"73812a70",
  1599 => x"81065152",
  1600 => x"71802e85",
  1601 => x"38728207",
  1602 => x"5372fc0c",
  1603 => x"865280e3",
  1604 => x"c4088338",
  1605 => x"845271ec",
  1606 => x"0cb1d804",
  1607 => x"800b80e3",
  1608 => x"c40c0290",
  1609 => x"050d0471",
  1610 => x"980c04ff",
  1611 => x"b00880e3",
  1612 => x"c40c0481",
  1613 => x"0bffb00c",
  1614 => x"04800bff",
  1615 => x"b00c0402",
  1616 => x"f4050db3",
  1617 => x"cd0480e3",
  1618 => x"c40881f0",
  1619 => x"2e098106",
  1620 => x"8a38810b",
  1621 => x"80e1f80c",
  1622 => x"b3cd0480",
  1623 => x"e3c40881",
  1624 => x"e02e0981",
  1625 => x"068a3881",
  1626 => x"0b80e1fc",
  1627 => x"0cb3cd04",
  1628 => x"80e3c408",
  1629 => x"5280e1fc",
  1630 => x"08802e89",
  1631 => x"3880e3c4",
  1632 => x"08818005",
  1633 => x"5271842c",
  1634 => x"728f0653",
  1635 => x"5380e1f8",
  1636 => x"08802e9a",
  1637 => x"38728429",
  1638 => x"80e1b805",
  1639 => x"72138171",
  1640 => x"2b700973",
  1641 => x"0806730c",
  1642 => x"515353b3",
  1643 => x"c1047284",
  1644 => x"2980e1b8",
  1645 => x"05721383",
  1646 => x"712b7208",
  1647 => x"07720c53",
  1648 => x"53800b80",
  1649 => x"e1fc0c80",
  1650 => x"0b80e1f8",
  1651 => x"0c80e3ec",
  1652 => x"51b4d42d",
  1653 => x"80e3c408",
  1654 => x"ff24feea",
  1655 => x"38800b80",
  1656 => x"e3c40c02",
  1657 => x"8c050d04",
  1658 => x"02f8050d",
  1659 => x"80e1b852",
  1660 => x"8f518072",
  1661 => x"70840554",
  1662 => x"0cff1151",
  1663 => x"708025f2",
  1664 => x"38028805",
  1665 => x"0d0402f0",
  1666 => x"050d7551",
  1667 => x"b2b92d70",
  1668 => x"822cfc06",
  1669 => x"80e1b811",
  1670 => x"72109e06",
  1671 => x"71087072",
  1672 => x"2a708306",
  1673 => x"82742b70",
  1674 => x"09740676",
  1675 => x"0c545156",
  1676 => x"57535153",
  1677 => x"b2b32d71",
  1678 => x"80e3c40c",
  1679 => x"0290050d",
  1680 => x"0402fc05",
  1681 => x"0d725180",
  1682 => x"710c800b",
  1683 => x"84120c02",
  1684 => x"84050d04",
  1685 => x"02f0050d",
  1686 => x"75700884",
  1687 => x"12085353",
  1688 => x"53ff5471",
  1689 => x"712ea838",
  1690 => x"b2b92d84",
  1691 => x"13087084",
  1692 => x"29148811",
  1693 => x"70087081",
  1694 => x"ff068418",
  1695 => x"08811187",
  1696 => x"06841a0c",
  1697 => x"53515551",
  1698 => x"5151b2b3",
  1699 => x"2d715473",
  1700 => x"80e3c40c",
  1701 => x"0290050d",
  1702 => x"0402f805",
  1703 => x"0db2b92d",
  1704 => x"e008708b",
  1705 => x"2a708106",
  1706 => x"51525270",
  1707 => x"802ea138",
  1708 => x"80e3ec08",
  1709 => x"70842980",
  1710 => x"e3f40573",
  1711 => x"81ff0671",
  1712 => x"0c515180",
  1713 => x"e3ec0881",
  1714 => x"11870680",
  1715 => x"e3ec0c51",
  1716 => x"800b80e4",
  1717 => x"940cb2ab",
  1718 => x"2db2b32d",
  1719 => x"0288050d",
  1720 => x"0402fc05",
  1721 => x"0db2b92d",
  1722 => x"810b80e4",
  1723 => x"940cb2b3",
  1724 => x"2d80e494",
  1725 => x"085170f9",
  1726 => x"38028405",
  1727 => x"0d0402fc",
  1728 => x"050d80e3",
  1729 => x"ec51b4c1",
  1730 => x"2db3e82d",
  1731 => x"b59951b2",
  1732 => x"a72d0284",
  1733 => x"050d0480",
  1734 => x"e4a00880",
  1735 => x"e3c40c04",
  1736 => x"02fc050d",
  1737 => x"810b80e2",
  1738 => x"840c8151",
  1739 => x"858d2d02",
  1740 => x"84050d04",
  1741 => x"02fc050d",
  1742 => x"b6be04b2",
  1743 => x"bf2d80f6",
  1744 => x"51b4862d",
  1745 => x"80e3c408",
  1746 => x"f23880da",
  1747 => x"51b4862d",
  1748 => x"80e3c408",
  1749 => x"e63880e3",
  1750 => x"c40880e2",
  1751 => x"840c80e3",
  1752 => x"c4085185",
  1753 => x"8d2d0284",
  1754 => x"050d0402",
  1755 => x"ec050d76",
  1756 => x"54805287",
  1757 => x"0b881580",
  1758 => x"f52d5653",
  1759 => x"74722483",
  1760 => x"38a05372",
  1761 => x"5183842d",
  1762 => x"81128b15",
  1763 => x"80f52d54",
  1764 => x"52727225",
  1765 => x"de380294",
  1766 => x"050d0402",
  1767 => x"f0050d80",
  1768 => x"e4a00854",
  1769 => x"81f92d80",
  1770 => x"0b80e4a4",
  1771 => x"0c730880",
  1772 => x"2e818938",
  1773 => x"820b80e3",
  1774 => x"d80c80e4",
  1775 => x"a4088f06",
  1776 => x"80e3d40c",
  1777 => x"73085271",
  1778 => x"832e9638",
  1779 => x"71832689",
  1780 => x"3871812e",
  1781 => x"b038b8a5",
  1782 => x"0471852e",
  1783 => x"a038b8a5",
  1784 => x"04881480",
  1785 => x"f52d8415",
  1786 => x"0880defc",
  1787 => x"53545286",
  1788 => x"a02d7184",
  1789 => x"29137008",
  1790 => x"5252b8a9",
  1791 => x"047351b6",
  1792 => x"eb2db8a5",
  1793 => x"0480e280",
  1794 => x"08881508",
  1795 => x"2c708106",
  1796 => x"51527180",
  1797 => x"2e883880",
  1798 => x"df8051b8",
  1799 => x"a20480df",
  1800 => x"845186a0",
  1801 => x"2d841408",
  1802 => x"5186a02d",
  1803 => x"80e4a408",
  1804 => x"810580e4",
  1805 => x"a40c8c14",
  1806 => x"54b7ad04",
  1807 => x"0290050d",
  1808 => x"047180e4",
  1809 => x"a00cb79b",
  1810 => x"2d80e4a4",
  1811 => x"08ff0580",
  1812 => x"e4a80c04",
  1813 => x"02e8050d",
  1814 => x"80e4a008",
  1815 => x"80e4ac08",
  1816 => x"575580f6",
  1817 => x"51b4862d",
  1818 => x"80e3c408",
  1819 => x"812a7081",
  1820 => x"06515271",
  1821 => x"802ea438",
  1822 => x"b8fe04b2",
  1823 => x"bf2d80f6",
  1824 => x"51b4862d",
  1825 => x"80e3c408",
  1826 => x"f23880e2",
  1827 => x"84088132",
  1828 => x"7080e284",
  1829 => x"0c705252",
  1830 => x"858d2d80",
  1831 => x"0b80e498",
  1832 => x"0c800b80",
  1833 => x"e49c0c80",
  1834 => x"e2840883",
  1835 => x"8e3880da",
  1836 => x"51b4862d",
  1837 => x"80e3c408",
  1838 => x"802e8c38",
  1839 => x"80e49808",
  1840 => x"81800780",
  1841 => x"e4980c80",
  1842 => x"d951b486",
  1843 => x"2d80e3c4",
  1844 => x"08802e8c",
  1845 => x"3880e498",
  1846 => x"0880c007",
  1847 => x"80e4980c",
  1848 => x"819451b4",
  1849 => x"862d80e3",
  1850 => x"c408802e",
  1851 => x"8b3880e4",
  1852 => x"98089007",
  1853 => x"80e4980c",
  1854 => x"819151b4",
  1855 => x"862d80e3",
  1856 => x"c408802e",
  1857 => x"8b3880e4",
  1858 => x"9808a007",
  1859 => x"80e4980c",
  1860 => x"81f551b4",
  1861 => x"862d80e3",
  1862 => x"c408802e",
  1863 => x"8b3880e4",
  1864 => x"98088107",
  1865 => x"80e4980c",
  1866 => x"81f251b4",
  1867 => x"862d80e3",
  1868 => x"c408802e",
  1869 => x"8b3880e4",
  1870 => x"98088207",
  1871 => x"80e4980c",
  1872 => x"81eb51b4",
  1873 => x"862d80e3",
  1874 => x"c408802e",
  1875 => x"8b3880e4",
  1876 => x"98088407",
  1877 => x"80e4980c",
  1878 => x"81f451b4",
  1879 => x"862d80e3",
  1880 => x"c408802e",
  1881 => x"8b3880e4",
  1882 => x"98088807",
  1883 => x"80e4980c",
  1884 => x"80d851b4",
  1885 => x"862d80e3",
  1886 => x"c408802e",
  1887 => x"8c3880e4",
  1888 => x"9c088180",
  1889 => x"0780e49c",
  1890 => x"0c9251b4",
  1891 => x"862d80e3",
  1892 => x"c408802e",
  1893 => x"8c3880e4",
  1894 => x"9c0880c0",
  1895 => x"0780e49c",
  1896 => x"0c9451b4",
  1897 => x"862d80e3",
  1898 => x"c408802e",
  1899 => x"8b3880e4",
  1900 => x"9c089007",
  1901 => x"80e49c0c",
  1902 => x"9151b486",
  1903 => x"2d80e3c4",
  1904 => x"08802e8b",
  1905 => x"3880e49c",
  1906 => x"08a00780",
  1907 => x"e49c0c9d",
  1908 => x"51b4862d",
  1909 => x"80e3c408",
  1910 => x"802e8b38",
  1911 => x"80e49c08",
  1912 => x"810780e4",
  1913 => x"9c0c9b51",
  1914 => x"b4862d80",
  1915 => x"e3c40880",
  1916 => x"2e8b3880",
  1917 => x"e49c0882",
  1918 => x"0780e49c",
  1919 => x"0c9c51b4",
  1920 => x"862d80e3",
  1921 => x"c408802e",
  1922 => x"8b3880e4",
  1923 => x"9c088407",
  1924 => x"80e49c0c",
  1925 => x"a351b486",
  1926 => x"2d80e3c4",
  1927 => x"08802e8b",
  1928 => x"3880e49c",
  1929 => x"08880780",
  1930 => x"e49c0c81",
  1931 => x"fd51b486",
  1932 => x"2d81fa51",
  1933 => x"b4862d80",
  1934 => x"c2960481",
  1935 => x"f551b486",
  1936 => x"2d80e3c4",
  1937 => x"08812a70",
  1938 => x"81065152",
  1939 => x"71802eb3",
  1940 => x"3880e4a8",
  1941 => x"08527180",
  1942 => x"2e8a38ff",
  1943 => x"1280e4a8",
  1944 => x"0cbd8304",
  1945 => x"80e4a408",
  1946 => x"1080e4a4",
  1947 => x"08057084",
  1948 => x"29165152",
  1949 => x"88120880",
  1950 => x"2e8938ff",
  1951 => x"51881208",
  1952 => x"52712d81",
  1953 => x"f251b486",
  1954 => x"2d80e3c4",
  1955 => x"08812a70",
  1956 => x"81065152",
  1957 => x"71802eb4",
  1958 => x"3880e4a4",
  1959 => x"08ff1180",
  1960 => x"e4a80856",
  1961 => x"53537372",
  1962 => x"258a3881",
  1963 => x"1480e4a8",
  1964 => x"0cbdcc04",
  1965 => x"72101370",
  1966 => x"84291651",
  1967 => x"52881208",
  1968 => x"802e8938",
  1969 => x"fe518812",
  1970 => x"0852712d",
  1971 => x"81fd51b4",
  1972 => x"862d80e3",
  1973 => x"c408812a",
  1974 => x"70810651",
  1975 => x"5271802e",
  1976 => x"b13880e4",
  1977 => x"a808802e",
  1978 => x"8a38800b",
  1979 => x"80e4a80c",
  1980 => x"be920480",
  1981 => x"e4a40810",
  1982 => x"80e4a408",
  1983 => x"05708429",
  1984 => x"16515288",
  1985 => x"1208802e",
  1986 => x"8938fd51",
  1987 => x"88120852",
  1988 => x"712d81fa",
  1989 => x"51b4862d",
  1990 => x"80e3c408",
  1991 => x"812a7081",
  1992 => x"06515271",
  1993 => x"802eb138",
  1994 => x"80e4a408",
  1995 => x"ff115452",
  1996 => x"80e4a808",
  1997 => x"73258938",
  1998 => x"7280e4a8",
  1999 => x"0cbed804",
  2000 => x"71101270",
  2001 => x"84291651",
  2002 => x"52881208",
  2003 => x"802e8938",
  2004 => x"fc518812",
  2005 => x"0852712d",
  2006 => x"80e4a808",
  2007 => x"70535473",
  2008 => x"802e8a38",
  2009 => x"8c15ff15",
  2010 => x"5555bedf",
  2011 => x"04820b80",
  2012 => x"e3d80c71",
  2013 => x"8f0680e3",
  2014 => x"d40c81eb",
  2015 => x"51b4862d",
  2016 => x"80e3c408",
  2017 => x"812a7081",
  2018 => x"06515271",
  2019 => x"802ead38",
  2020 => x"7408852e",
  2021 => x"098106a4",
  2022 => x"38881580",
  2023 => x"f52dff05",
  2024 => x"52718816",
  2025 => x"81b72d71",
  2026 => x"982b5271",
  2027 => x"80258838",
  2028 => x"800b8816",
  2029 => x"81b72d74",
  2030 => x"51b6eb2d",
  2031 => x"81f451b4",
  2032 => x"862d80e3",
  2033 => x"c408812a",
  2034 => x"70810651",
  2035 => x"5271802e",
  2036 => x"b3387408",
  2037 => x"852e0981",
  2038 => x"06aa3888",
  2039 => x"1580f52d",
  2040 => x"81055271",
  2041 => x"881681b7",
  2042 => x"2d7181ff",
  2043 => x"068b1680",
  2044 => x"f52d5452",
  2045 => x"72722787",
  2046 => x"38728816",
  2047 => x"81b72d74",
  2048 => x"51b6eb2d",
  2049 => x"80da51b4",
  2050 => x"862d80e3",
  2051 => x"c408812a",
  2052 => x"70810651",
  2053 => x"5271802e",
  2054 => x"81b33880",
  2055 => x"e4a00880",
  2056 => x"e4a80855",
  2057 => x"5373802e",
  2058 => x"8b388c13",
  2059 => x"ff155553",
  2060 => x"80c0a504",
  2061 => x"72085271",
  2062 => x"822ea838",
  2063 => x"7182268a",
  2064 => x"3871812e",
  2065 => x"ad3880c1",
  2066 => x"cd047183",
  2067 => x"2eb73871",
  2068 => x"842e0981",
  2069 => x"0680f638",
  2070 => x"88130851",
  2071 => x"b8c12d80",
  2072 => x"c1cd0480",
  2073 => x"e4a80851",
  2074 => x"88130852",
  2075 => x"712d80c1",
  2076 => x"cd04810b",
  2077 => x"8814082b",
  2078 => x"80e28008",
  2079 => x"3280e280",
  2080 => x"0c80c1a0",
  2081 => x"04881380",
  2082 => x"f52d8105",
  2083 => x"8b1480f5",
  2084 => x"2d535471",
  2085 => x"74248338",
  2086 => x"80547388",
  2087 => x"1481b72d",
  2088 => x"b79b2d80",
  2089 => x"c1cd0475",
  2090 => x"08802ea4",
  2091 => x"38750851",
  2092 => x"b4862d80",
  2093 => x"e3c40881",
  2094 => x"06527180",
  2095 => x"2e8c3880",
  2096 => x"e4a80851",
  2097 => x"84160852",
  2098 => x"712d8816",
  2099 => x"5675d838",
  2100 => x"8054800b",
  2101 => x"80e3d80c",
  2102 => x"738f0680",
  2103 => x"e3d40ca0",
  2104 => x"527380e4",
  2105 => x"a8082e09",
  2106 => x"81069938",
  2107 => x"80e4a408",
  2108 => x"ff057432",
  2109 => x"70098105",
  2110 => x"7072079f",
  2111 => x"2a917131",
  2112 => x"51515353",
  2113 => x"71518384",
  2114 => x"2d811454",
  2115 => x"8e7425c2",
  2116 => x"3880e284",
  2117 => x"08527180",
  2118 => x"e3c40c02",
  2119 => x"98050d04",
  2120 => x"02f4050d",
  2121 => x"d45281ff",
  2122 => x"720c7108",
  2123 => x"5381ff72",
  2124 => x"0c72882b",
  2125 => x"83fe8006",
  2126 => x"72087081",
  2127 => x"ff065152",
  2128 => x"5381ff72",
  2129 => x"0c727107",
  2130 => x"882b7208",
  2131 => x"7081ff06",
  2132 => x"51525381",
  2133 => x"ff720c72",
  2134 => x"7107882b",
  2135 => x"72087081",
  2136 => x"ff067207",
  2137 => x"80e3c40c",
  2138 => x"5253028c",
  2139 => x"050d0402",
  2140 => x"f4050d74",
  2141 => x"767181ff",
  2142 => x"06d40c53",
  2143 => x"5380e4b0",
  2144 => x"08853871",
  2145 => x"892b5271",
  2146 => x"982ad40c",
  2147 => x"71902a70",
  2148 => x"81ff06d4",
  2149 => x"0c517188",
  2150 => x"2a7081ff",
  2151 => x"06d40c51",
  2152 => x"7181ff06",
  2153 => x"d40c7290",
  2154 => x"2a7081ff",
  2155 => x"06d40c51",
  2156 => x"d4087081",
  2157 => x"ff065151",
  2158 => x"82b8bf52",
  2159 => x"7081ff2e",
  2160 => x"09810694",
  2161 => x"3881ff0b",
  2162 => x"d40cd408",
  2163 => x"7081ff06",
  2164 => x"ff145451",
  2165 => x"5171e538",
  2166 => x"7080e3c4",
  2167 => x"0c028c05",
  2168 => x"0d0402fc",
  2169 => x"050d81c7",
  2170 => x"5181ff0b",
  2171 => x"d40cff11",
  2172 => x"51708025",
  2173 => x"f4380284",
  2174 => x"050d0402",
  2175 => x"f4050d81",
  2176 => x"ff0bd40c",
  2177 => x"93538052",
  2178 => x"87fc80c1",
  2179 => x"5180c2ef",
  2180 => x"2d80e3c4",
  2181 => x"088c3881",
  2182 => x"ff0bd40c",
  2183 => x"815380c4",
  2184 => x"ac0480c3",
  2185 => x"e22dff13",
  2186 => x"5372db38",
  2187 => x"7280e3c4",
  2188 => x"0c028c05",
  2189 => x"0d0402ec",
  2190 => x"050d810b",
  2191 => x"80e4b00c",
  2192 => x"8454d008",
  2193 => x"708f2a70",
  2194 => x"81065151",
  2195 => x"5372f338",
  2196 => x"72d00c80",
  2197 => x"c3e22d80",
  2198 => x"df885186",
  2199 => x"a02dd008",
  2200 => x"708f2a70",
  2201 => x"81065151",
  2202 => x"5372f338",
  2203 => x"810bd00c",
  2204 => x"b1538052",
  2205 => x"84d480c0",
  2206 => x"5180c2ef",
  2207 => x"2d80e3c4",
  2208 => x"08812e94",
  2209 => x"3872822e",
  2210 => x"80c438ff",
  2211 => x"135372e2",
  2212 => x"38ff1454",
  2213 => x"73ffab38",
  2214 => x"80c3e22d",
  2215 => x"83aa5284",
  2216 => x"9c80c851",
  2217 => x"80c2ef2d",
  2218 => x"80e3c408",
  2219 => x"812e0981",
  2220 => x"06943880",
  2221 => x"c2a02d80",
  2222 => x"e3c40883",
  2223 => x"ffff0653",
  2224 => x"7283aa2e",
  2225 => x"a33880c3",
  2226 => x"fb2d80c5",
  2227 => x"e20480df",
  2228 => x"945186a0",
  2229 => x"2d805380",
  2230 => x"c7c00480",
  2231 => x"dfac5186",
  2232 => x"a02d8054",
  2233 => x"80c79004",
  2234 => x"81ff0bd4",
  2235 => x"0cb15480",
  2236 => x"c3e22d8f",
  2237 => x"cf538052",
  2238 => x"87fc80f7",
  2239 => x"5180c2ef",
  2240 => x"2d80e3c4",
  2241 => x"085580e3",
  2242 => x"c408812e",
  2243 => x"0981069e",
  2244 => x"3881ff0b",
  2245 => x"d40c820a",
  2246 => x"52849c80",
  2247 => x"e95180c2",
  2248 => x"ef2d80e3",
  2249 => x"c408802e",
  2250 => x"8f3880c3",
  2251 => x"e22dff13",
  2252 => x"5372c338",
  2253 => x"80c78304",
  2254 => x"81ff0bd4",
  2255 => x"0c80e3c4",
  2256 => x"085287fc",
  2257 => x"80fa5180",
  2258 => x"c2ef2d80",
  2259 => x"e3c408b3",
  2260 => x"3881ff0b",
  2261 => x"d40cd408",
  2262 => x"5381ff0b",
  2263 => x"d40c81ff",
  2264 => x"0bd40c81",
  2265 => x"ff0bd40c",
  2266 => x"81ff0bd4",
  2267 => x"0c72862a",
  2268 => x"70810676",
  2269 => x"56515372",
  2270 => x"973880e3",
  2271 => x"c4085480",
  2272 => x"c7900473",
  2273 => x"822efed3",
  2274 => x"38ff1454",
  2275 => x"73fee038",
  2276 => x"7380e4b0",
  2277 => x"0c738c38",
  2278 => x"815287fc",
  2279 => x"80d05180",
  2280 => x"c2ef2d81",
  2281 => x"ff0bd40c",
  2282 => x"d008708f",
  2283 => x"2a708106",
  2284 => x"51515372",
  2285 => x"f33872d0",
  2286 => x"0c81ff0b",
  2287 => x"d40c8153",
  2288 => x"7280e3c4",
  2289 => x"0c029405",
  2290 => x"0d0402e8",
  2291 => x"050d7855",
  2292 => x"805681ff",
  2293 => x"0bd40cd0",
  2294 => x"08708f2a",
  2295 => x"70810651",
  2296 => x"515372f3",
  2297 => x"3882810b",
  2298 => x"d00c81ff",
  2299 => x"0bd40c77",
  2300 => x"5287fc80",
  2301 => x"d15180c2",
  2302 => x"ef2d80db",
  2303 => x"c6df5480",
  2304 => x"e3c40880",
  2305 => x"2e8c3880",
  2306 => x"dfcc5186",
  2307 => x"a02d80c8",
  2308 => x"e80481ff",
  2309 => x"0bd40cd4",
  2310 => x"087081ff",
  2311 => x"06515372",
  2312 => x"81fe2e09",
  2313 => x"8106a038",
  2314 => x"80ff5380",
  2315 => x"c2a02d80",
  2316 => x"e3c40875",
  2317 => x"70840557",
  2318 => x"0cff1353",
  2319 => x"728025eb",
  2320 => x"38815680",
  2321 => x"c8cd04ff",
  2322 => x"145473c6",
  2323 => x"3881ff0b",
  2324 => x"d40c81ff",
  2325 => x"0bd40cd0",
  2326 => x"08708f2a",
  2327 => x"70810651",
  2328 => x"515372f3",
  2329 => x"3872d00c",
  2330 => x"7580e3c4",
  2331 => x"0c029805",
  2332 => x"0d0402e8",
  2333 => x"050d7779",
  2334 => x"7b585555",
  2335 => x"80537276",
  2336 => x"25a53874",
  2337 => x"70810556",
  2338 => x"80f52d74",
  2339 => x"70810556",
  2340 => x"80f52d52",
  2341 => x"5271712e",
  2342 => x"87388151",
  2343 => x"80c9a904",
  2344 => x"81135380",
  2345 => x"c8fe0480",
  2346 => x"517080e3",
  2347 => x"c40c0298",
  2348 => x"050d0402",
  2349 => x"ec050d76",
  2350 => x"5574802e",
  2351 => x"80c4389a",
  2352 => x"1580e02d",
  2353 => x"5180d7ee",
  2354 => x"2d80e3c4",
  2355 => x"0880e3c4",
  2356 => x"0880eae4",
  2357 => x"0c80e3c4",
  2358 => x"08545480",
  2359 => x"eac00880",
  2360 => x"2e9b3894",
  2361 => x"1580e02d",
  2362 => x"5180d7ee",
  2363 => x"2d80e3c4",
  2364 => x"08902b83",
  2365 => x"fff00a06",
  2366 => x"70750751",
  2367 => x"537280ea",
  2368 => x"e40c80ea",
  2369 => x"e4085372",
  2370 => x"802e9e38",
  2371 => x"80eab808",
  2372 => x"fe147129",
  2373 => x"80eacc08",
  2374 => x"0580eae8",
  2375 => x"0c70842b",
  2376 => x"80eac40c",
  2377 => x"5480cad8",
  2378 => x"0480ead0",
  2379 => x"0880eae4",
  2380 => x"0c80ead4",
  2381 => x"0880eae8",
  2382 => x"0c80eac0",
  2383 => x"08802e8c",
  2384 => x"3880eab8",
  2385 => x"08842b53",
  2386 => x"80cad304",
  2387 => x"80ead808",
  2388 => x"842b5372",
  2389 => x"80eac40c",
  2390 => x"0294050d",
  2391 => x"0402d805",
  2392 => x"0d800b80",
  2393 => x"eac00c84",
  2394 => x"5480c4b6",
  2395 => x"2d80e3c4",
  2396 => x"08802e99",
  2397 => x"3880e4b4",
  2398 => x"52805180",
  2399 => x"c7ca2d80",
  2400 => x"e3c40880",
  2401 => x"2e8738fe",
  2402 => x"5480cb95",
  2403 => x"04ff1454",
  2404 => x"738024d5",
  2405 => x"38738e38",
  2406 => x"80dfdc51",
  2407 => x"86a02d73",
  2408 => x"5580d0f9",
  2409 => x"04805681",
  2410 => x"0b80eaec",
  2411 => x"0c885380",
  2412 => x"dff05280",
  2413 => x"e4ea5180",
  2414 => x"c8f22d80",
  2415 => x"e3c40876",
  2416 => x"2e098106",
  2417 => x"893880e3",
  2418 => x"c40880ea",
  2419 => x"ec0c8853",
  2420 => x"80dffc52",
  2421 => x"80e58651",
  2422 => x"80c8f22d",
  2423 => x"80e3c408",
  2424 => x"893880e3",
  2425 => x"c40880ea",
  2426 => x"ec0c80ea",
  2427 => x"ec08802e",
  2428 => x"81853880",
  2429 => x"e7fa0b80",
  2430 => x"f52d80e7",
  2431 => x"fb0b80f5",
  2432 => x"2d71982b",
  2433 => x"71902b07",
  2434 => x"80e7fc0b",
  2435 => x"80f52d70",
  2436 => x"882b7207",
  2437 => x"80e7fd0b",
  2438 => x"80f52d71",
  2439 => x"0780e8b2",
  2440 => x"0b80f52d",
  2441 => x"80e8b30b",
  2442 => x"80f52d71",
  2443 => x"882b0753",
  2444 => x"5f54525a",
  2445 => x"56575573",
  2446 => x"81abaa2e",
  2447 => x"09810690",
  2448 => x"38755180",
  2449 => x"d7bd2d80",
  2450 => x"e3c40856",
  2451 => x"80ccdf04",
  2452 => x"7382d4d5",
  2453 => x"2e893880",
  2454 => x"e0885180",
  2455 => x"cdaf0480",
  2456 => x"e4b45275",
  2457 => x"5180c7ca",
  2458 => x"2d80e3c4",
  2459 => x"085580e3",
  2460 => x"c408802e",
  2461 => x"84833888",
  2462 => x"5380dffc",
  2463 => x"5280e586",
  2464 => x"5180c8f2",
  2465 => x"2d80e3c4",
  2466 => x"088b3881",
  2467 => x"0b80eac0",
  2468 => x"0c80cdb6",
  2469 => x"04885380",
  2470 => x"dff05280",
  2471 => x"e4ea5180",
  2472 => x"c8f22d80",
  2473 => x"e3c40880",
  2474 => x"2e8c3880",
  2475 => x"e09c5186",
  2476 => x"a02d80ce",
  2477 => x"950480e8",
  2478 => x"b20b80f5",
  2479 => x"2d547380",
  2480 => x"d52e0981",
  2481 => x"0680ce38",
  2482 => x"80e8b30b",
  2483 => x"80f52d54",
  2484 => x"7381aa2e",
  2485 => x"098106bd",
  2486 => x"38800b80",
  2487 => x"e4b40b80",
  2488 => x"f52d5654",
  2489 => x"7481e92e",
  2490 => x"83388154",
  2491 => x"7481eb2e",
  2492 => x"8c388055",
  2493 => x"73752e09",
  2494 => x"810682fd",
  2495 => x"3880e4bf",
  2496 => x"0b80f52d",
  2497 => x"55748e38",
  2498 => x"80e4c00b",
  2499 => x"80f52d54",
  2500 => x"73822e87",
  2501 => x"38805580",
  2502 => x"d0f90480",
  2503 => x"e4c10b80",
  2504 => x"f52d7080",
  2505 => x"eab80cff",
  2506 => x"0580eabc",
  2507 => x"0c80e4c2",
  2508 => x"0b80f52d",
  2509 => x"80e4c30b",
  2510 => x"80f52d58",
  2511 => x"76057782",
  2512 => x"80290570",
  2513 => x"80eac80c",
  2514 => x"80e4c40b",
  2515 => x"80f52d70",
  2516 => x"80eadc0c",
  2517 => x"80eac008",
  2518 => x"59575876",
  2519 => x"802e81b9",
  2520 => x"38885380",
  2521 => x"dffc5280",
  2522 => x"e5865180",
  2523 => x"c8f22d80",
  2524 => x"e3c40882",
  2525 => x"843880ea",
  2526 => x"b8087084",
  2527 => x"2b80eac4",
  2528 => x"0c7080ea",
  2529 => x"d80c80e4",
  2530 => x"d90b80f5",
  2531 => x"2d80e4d8",
  2532 => x"0b80f52d",
  2533 => x"71828029",
  2534 => x"0580e4da",
  2535 => x"0b80f52d",
  2536 => x"70848080",
  2537 => x"291280e4",
  2538 => x"db0b80f5",
  2539 => x"2d708180",
  2540 => x"0a291270",
  2541 => x"80eae00c",
  2542 => x"80eadc08",
  2543 => x"712980ea",
  2544 => x"c8080570",
  2545 => x"80eacc0c",
  2546 => x"80e4e10b",
  2547 => x"80f52d80",
  2548 => x"e4e00b80",
  2549 => x"f52d7182",
  2550 => x"80290580",
  2551 => x"e4e20b80",
  2552 => x"f52d7084",
  2553 => x"80802912",
  2554 => x"80e4e30b",
  2555 => x"80f52d70",
  2556 => x"982b81f0",
  2557 => x"0a067205",
  2558 => x"7080ead0",
  2559 => x"0cfe117e",
  2560 => x"29770580",
  2561 => x"ead40c52",
  2562 => x"59524354",
  2563 => x"5e515259",
  2564 => x"525d5759",
  2565 => x"5780d0f1",
  2566 => x"0480e4c6",
  2567 => x"0b80f52d",
  2568 => x"80e4c50b",
  2569 => x"80f52d71",
  2570 => x"82802905",
  2571 => x"7080eac4",
  2572 => x"0c70a029",
  2573 => x"83ff0570",
  2574 => x"892a7080",
  2575 => x"ead80c80",
  2576 => x"e4cb0b80",
  2577 => x"f52d80e4",
  2578 => x"ca0b80f5",
  2579 => x"2d718280",
  2580 => x"29057080",
  2581 => x"eae00c7b",
  2582 => x"71291e70",
  2583 => x"80ead40c",
  2584 => x"7d80ead0",
  2585 => x"0c730580",
  2586 => x"eacc0c55",
  2587 => x"5e515155",
  2588 => x"55805180",
  2589 => x"c9b32d81",
  2590 => x"557480e3",
  2591 => x"c40c02a8",
  2592 => x"050d0402",
  2593 => x"ec050d76",
  2594 => x"70872c71",
  2595 => x"80ff0655",
  2596 => x"565480ea",
  2597 => x"c0088a38",
  2598 => x"73882c74",
  2599 => x"81ff0654",
  2600 => x"5580e4b4",
  2601 => x"5280eac8",
  2602 => x"08155180",
  2603 => x"c7ca2d80",
  2604 => x"e3c40854",
  2605 => x"80e3c408",
  2606 => x"802ebb38",
  2607 => x"80eac008",
  2608 => x"802e9c38",
  2609 => x"72842980",
  2610 => x"e4b40570",
  2611 => x"08525380",
  2612 => x"d7bd2d80",
  2613 => x"e3c408f0",
  2614 => x"0a065380",
  2615 => x"d1f40472",
  2616 => x"1080e4b4",
  2617 => x"057080e0",
  2618 => x"2d525380",
  2619 => x"d7ee2d80",
  2620 => x"e3c40853",
  2621 => x"72547380",
  2622 => x"e3c40c02",
  2623 => x"94050d04",
  2624 => x"02e0050d",
  2625 => x"7970842c",
  2626 => x"80eae808",
  2627 => x"05718f06",
  2628 => x"52555372",
  2629 => x"8b3880e4",
  2630 => x"b4527351",
  2631 => x"80c7ca2d",
  2632 => x"72a02980",
  2633 => x"e4b40554",
  2634 => x"807480f5",
  2635 => x"2d565374",
  2636 => x"732e8338",
  2637 => x"81537481",
  2638 => x"e52e81f5",
  2639 => x"38817074",
  2640 => x"06545872",
  2641 => x"802e81e9",
  2642 => x"388b1480",
  2643 => x"f52d7083",
  2644 => x"2a790658",
  2645 => x"56769c38",
  2646 => x"80e28808",
  2647 => x"53728938",
  2648 => x"7280e8b4",
  2649 => x"0b81b72d",
  2650 => x"7680e288",
  2651 => x"0c735380",
  2652 => x"d4b30475",
  2653 => x"8f2e0981",
  2654 => x"0681b638",
  2655 => x"749f068d",
  2656 => x"2980e8a7",
  2657 => x"11515381",
  2658 => x"1480f52d",
  2659 => x"73708105",
  2660 => x"5581b72d",
  2661 => x"831480f5",
  2662 => x"2d737081",
  2663 => x"055581b7",
  2664 => x"2d851480",
  2665 => x"f52d7370",
  2666 => x"81055581",
  2667 => x"b72d8714",
  2668 => x"80f52d73",
  2669 => x"70810555",
  2670 => x"81b72d89",
  2671 => x"1480f52d",
  2672 => x"73708105",
  2673 => x"5581b72d",
  2674 => x"8e1480f5",
  2675 => x"2d737081",
  2676 => x"055581b7",
  2677 => x"2d901480",
  2678 => x"f52d7370",
  2679 => x"81055581",
  2680 => x"b72d9214",
  2681 => x"80f52d73",
  2682 => x"70810555",
  2683 => x"81b72d94",
  2684 => x"1480f52d",
  2685 => x"73708105",
  2686 => x"5581b72d",
  2687 => x"961480f5",
  2688 => x"2d737081",
  2689 => x"055581b7",
  2690 => x"2d981480",
  2691 => x"f52d7370",
  2692 => x"81055581",
  2693 => x"b72d9c14",
  2694 => x"80f52d73",
  2695 => x"70810555",
  2696 => x"81b72d9e",
  2697 => x"1480f52d",
  2698 => x"7381b72d",
  2699 => x"7780e288",
  2700 => x"0c805372",
  2701 => x"80e3c40c",
  2702 => x"02a0050d",
  2703 => x"0402cc05",
  2704 => x"0d7e605e",
  2705 => x"5a800b80",
  2706 => x"eae40880",
  2707 => x"eae80859",
  2708 => x"5c568058",
  2709 => x"80eac408",
  2710 => x"782e81be",
  2711 => x"38778f06",
  2712 => x"a0175754",
  2713 => x"73923880",
  2714 => x"e4b45276",
  2715 => x"51811757",
  2716 => x"80c7ca2d",
  2717 => x"80e4b456",
  2718 => x"807680f5",
  2719 => x"2d565474",
  2720 => x"742e8338",
  2721 => x"81547481",
  2722 => x"e52e8182",
  2723 => x"38817075",
  2724 => x"06555c73",
  2725 => x"802e80f6",
  2726 => x"388b1680",
  2727 => x"f52d9806",
  2728 => x"597880ea",
  2729 => x"388b537c",
  2730 => x"52755180",
  2731 => x"c8f22d80",
  2732 => x"e3c40880",
  2733 => x"d9389c16",
  2734 => x"085180d7",
  2735 => x"bd2d80e3",
  2736 => x"c408841b",
  2737 => x"0c9a1680",
  2738 => x"e02d5180",
  2739 => x"d7ee2d80",
  2740 => x"e3c40880",
  2741 => x"e3c40888",
  2742 => x"1c0c80e3",
  2743 => x"c4085555",
  2744 => x"80eac008",
  2745 => x"802e9a38",
  2746 => x"941680e0",
  2747 => x"2d5180d7",
  2748 => x"ee2d80e3",
  2749 => x"c408902b",
  2750 => x"83fff00a",
  2751 => x"06701651",
  2752 => x"5473881b",
  2753 => x"0c787a0c",
  2754 => x"7b5480d6",
  2755 => x"d8048118",
  2756 => x"5880eac4",
  2757 => x"087826fe",
  2758 => x"c43880ea",
  2759 => x"c008802e",
  2760 => x"b5387a51",
  2761 => x"80d1832d",
  2762 => x"80e3c408",
  2763 => x"80e3c408",
  2764 => x"80ffffff",
  2765 => x"f806555b",
  2766 => x"7380ffff",
  2767 => x"fff82e96",
  2768 => x"3880e3c4",
  2769 => x"08fe0580",
  2770 => x"eab80829",
  2771 => x"80eacc08",
  2772 => x"055780d4",
  2773 => x"d2048054",
  2774 => x"7380e3c4",
  2775 => x"0c02b405",
  2776 => x"0d0402f4",
  2777 => x"050d7470",
  2778 => x"08810571",
  2779 => x"0c700880",
  2780 => x"eabc0806",
  2781 => x"53537190",
  2782 => x"38881308",
  2783 => x"5180d183",
  2784 => x"2d80e3c4",
  2785 => x"0888140c",
  2786 => x"810b80e3",
  2787 => x"c40c028c",
  2788 => x"050d0402",
  2789 => x"f0050d75",
  2790 => x"881108fe",
  2791 => x"0580eab8",
  2792 => x"082980ea",
  2793 => x"cc081172",
  2794 => x"0880eabc",
  2795 => x"08060579",
  2796 => x"55535454",
  2797 => x"80c7ca2d",
  2798 => x"0290050d",
  2799 => x"0402f405",
  2800 => x"0d747088",
  2801 => x"2a83fe80",
  2802 => x"06707298",
  2803 => x"2a077288",
  2804 => x"2b87fc80",
  2805 => x"80067398",
  2806 => x"2b81f00a",
  2807 => x"06717307",
  2808 => x"0780e3c4",
  2809 => x"0c565153",
  2810 => x"51028c05",
  2811 => x"0d0402f8",
  2812 => x"050d028e",
  2813 => x"0580f52d",
  2814 => x"74882b07",
  2815 => x"7083ffff",
  2816 => x"0680e3c4",
  2817 => x"0c510288",
  2818 => x"050d0402",
  2819 => x"f4050d74",
  2820 => x"76785354",
  2821 => x"52807125",
  2822 => x"97387270",
  2823 => x"81055480",
  2824 => x"f52d7270",
  2825 => x"81055481",
  2826 => x"b72dff11",
  2827 => x"5170eb38",
  2828 => x"807281b7",
  2829 => x"2d028c05",
  2830 => x"0d0402e8",
  2831 => x"050d7756",
  2832 => x"80705654",
  2833 => x"737624b7",
  2834 => x"3880eac4",
  2835 => x"08742eaf",
  2836 => x"38735180",
  2837 => x"d2802d80",
  2838 => x"e3c40880",
  2839 => x"e3c40809",
  2840 => x"81057080",
  2841 => x"e3c40807",
  2842 => x"9f2a7705",
  2843 => x"81175757",
  2844 => x"53537476",
  2845 => x"24893880",
  2846 => x"eac40874",
  2847 => x"26d33872",
  2848 => x"80e3c40c",
  2849 => x"0298050d",
  2850 => x"0402f005",
  2851 => x"0d80e3c0",
  2852 => x"08165180",
  2853 => x"d8ba2d80",
  2854 => x"e3c40880",
  2855 => x"2ea0388b",
  2856 => x"5380e3c4",
  2857 => x"085280e8",
  2858 => x"b45180d8",
  2859 => x"8b2d80ea",
  2860 => x"f0085473",
  2861 => x"802e8738",
  2862 => x"80e8b451",
  2863 => x"732d0290",
  2864 => x"050d0402",
  2865 => x"dc050d80",
  2866 => x"705a5574",
  2867 => x"80e3c008",
  2868 => x"25b53880",
  2869 => x"eac40875",
  2870 => x"2ead3878",
  2871 => x"5180d280",
  2872 => x"2d80e3c4",
  2873 => x"08098105",
  2874 => x"7080e3c4",
  2875 => x"08079f2a",
  2876 => x"7605811b",
  2877 => x"5b565474",
  2878 => x"80e3c008",
  2879 => x"25893880",
  2880 => x"eac40879",
  2881 => x"26d53880",
  2882 => x"557880ea",
  2883 => x"c4082781",
  2884 => x"e4387851",
  2885 => x"80d2802d",
  2886 => x"80e3c408",
  2887 => x"802e81b4",
  2888 => x"3880e3c4",
  2889 => x"088b0580",
  2890 => x"f52d7084",
  2891 => x"2a708106",
  2892 => x"77107884",
  2893 => x"2b80e8b4",
  2894 => x"0b80f52d",
  2895 => x"5c5c5351",
  2896 => x"55567380",
  2897 => x"2e80ce38",
  2898 => x"7416822b",
  2899 => x"80dc990b",
  2900 => x"80e29412",
  2901 => x"0c547775",
  2902 => x"311080ea",
  2903 => x"f4115556",
  2904 => x"90747081",
  2905 => x"055681b7",
  2906 => x"2da07481",
  2907 => x"b72d7681",
  2908 => x"ff068116",
  2909 => x"58547380",
  2910 => x"2e8b389c",
  2911 => x"5380e8b4",
  2912 => x"5280db8c",
  2913 => x"048b5380",
  2914 => x"e3c40852",
  2915 => x"80eaf616",
  2916 => x"5180dbca",
  2917 => x"04741682",
  2918 => x"2b80d989",
  2919 => x"0b80e294",
  2920 => x"120c5476",
  2921 => x"81ff0681",
  2922 => x"16585473",
  2923 => x"802e8b38",
  2924 => x"9c5380e8",
  2925 => x"b45280db",
  2926 => x"c1048b53",
  2927 => x"80e3c408",
  2928 => x"52777531",
  2929 => x"1080eaf4",
  2930 => x"05517655",
  2931 => x"80d88b2d",
  2932 => x"80dbe904",
  2933 => x"74902975",
  2934 => x"31701080",
  2935 => x"eaf40551",
  2936 => x"5480e3c4",
  2937 => x"087481b7",
  2938 => x"2d811959",
  2939 => x"748b24a4",
  2940 => x"3880da89",
  2941 => x"04749029",
  2942 => x"75317010",
  2943 => x"80eaf405",
  2944 => x"8c773157",
  2945 => x"51548074",
  2946 => x"81b72d9e",
  2947 => x"14ff1656",
  2948 => x"5474f338",
  2949 => x"02a4050d",
  2950 => x"0402fc05",
  2951 => x"0d80e3c0",
  2952 => x"08135180",
  2953 => x"d8ba2d80",
  2954 => x"e3c40880",
  2955 => x"2e8a3880",
  2956 => x"e3c40851",
  2957 => x"80c9b32d",
  2958 => x"800b80e3",
  2959 => x"c00c80d9",
  2960 => x"c32db79b",
  2961 => x"2d028405",
  2962 => x"0d0402fc",
  2963 => x"050d7251",
  2964 => x"70fd2eb2",
  2965 => x"3870fd24",
  2966 => x"8b3870fc",
  2967 => x"2e80d038",
  2968 => x"80ddb904",
  2969 => x"70fe2eb9",
  2970 => x"3870ff2e",
  2971 => x"09810680",
  2972 => x"c83880e3",
  2973 => x"c0085170",
  2974 => x"802ebe38",
  2975 => x"ff1180e3",
  2976 => x"c00c80dd",
  2977 => x"b90480e3",
  2978 => x"c008f005",
  2979 => x"7080e3c0",
  2980 => x"0c517080",
  2981 => x"25a33880",
  2982 => x"0b80e3c0",
  2983 => x"0c80ddb9",
  2984 => x"0480e3c0",
  2985 => x"08810580",
  2986 => x"e3c00c80",
  2987 => x"ddb90480",
  2988 => x"e3c00890",
  2989 => x"0580e3c0",
  2990 => x"0c80d9c3",
  2991 => x"2db79b2d",
  2992 => x"0284050d",
  2993 => x"0402fc05",
  2994 => x"0d800b80",
  2995 => x"e3c00c80",
  2996 => x"d9c32db6",
  2997 => x"972d80e3",
  2998 => x"c40880e3",
  2999 => x"b00c80e2",
  3000 => x"8c51b8c1",
  3001 => x"2d028405",
  3002 => x"0d047180",
  3003 => x"eaf00c04",
  3004 => x"00ffffff",
  3005 => x"ff00ffff",
  3006 => x"ffff00ff",
  3007 => x"ffffff00",
  3008 => x"52657365",
  3009 => x"74000000",
  3010 => x"5363616e",
  3011 => x"6c696e65",
  3012 => x"73000000",
  3013 => x"48513258",
  3014 => x"2046696c",
  3015 => x"74657200",
  3016 => x"50312053",
  3017 => x"656c6563",
  3018 => x"74000000",
  3019 => x"50312053",
  3020 => x"74617274",
  3021 => x"00000000",
  3022 => x"4c6f6164",
  3023 => x"20524f4d",
  3024 => x"20100000",
  3025 => x"45786974",
  3026 => x"00000000",
  3027 => x"524f4d20",
  3028 => x"6c6f6164",
  3029 => x"696e6720",
  3030 => x"6661696c",
  3031 => x"65640000",
  3032 => x"4f4b0000",
  3033 => x"496e6974",
  3034 => x"69616c69",
  3035 => x"7a696e67",
  3036 => x"20534420",
  3037 => x"63617264",
  3038 => x"0a000000",
  3039 => x"16200000",
  3040 => x"14200000",
  3041 => x"15200000",
  3042 => x"53442069",
  3043 => x"6e69742e",
  3044 => x"2e2e0a00",
  3045 => x"53442063",
  3046 => x"61726420",
  3047 => x"72657365",
  3048 => x"74206661",
  3049 => x"696c6564",
  3050 => x"210a0000",
  3051 => x"53444843",
  3052 => x"20657272",
  3053 => x"6f72210a",
  3054 => x"00000000",
  3055 => x"57726974",
  3056 => x"65206661",
  3057 => x"696c6564",
  3058 => x"0a000000",
  3059 => x"52656164",
  3060 => x"20666169",
  3061 => x"6c65640a",
  3062 => x"00000000",
  3063 => x"43617264",
  3064 => x"20696e69",
  3065 => x"74206661",
  3066 => x"696c6564",
  3067 => x"0a000000",
  3068 => x"46415431",
  3069 => x"36202020",
  3070 => x"00000000",
  3071 => x"46415433",
  3072 => x"32202020",
  3073 => x"00000000",
  3074 => x"4e6f2070",
  3075 => x"61727469",
  3076 => x"74696f6e",
  3077 => x"20736967",
  3078 => x"0a000000",
  3079 => x"42616420",
  3080 => x"70617274",
  3081 => x"0a000000",
  3082 => x"4261636b",
  3083 => x"00000000",
  3084 => x"00000002",
  3085 => x"00000002",
  3086 => x"00002f00",
  3087 => x"0000035a",
  3088 => x"00000001",
  3089 => x"00002f08",
  3090 => x"00000000",
  3091 => x"00000001",
  3092 => x"00002f14",
  3093 => x"00000001",
  3094 => x"00000002",
  3095 => x"00002f20",
  3096 => x"0000036e",
  3097 => x"00000002",
  3098 => x"00002f2c",
  3099 => x"00000a3f",
  3100 => x"00000002",
  3101 => x"00002f38",
  3102 => x"00002ec5",
  3103 => x"00000002",
  3104 => x"00002f44",
  3105 => x"00001b34",
  3106 => x"00000000",
  3107 => x"00000000",
  3108 => x"00000000",
  3109 => x"00000004",
  3110 => x"00002f4c",
  3111 => x"00003094",
  3112 => x"00000004",
  3113 => x"00002f60",
  3114 => x"00003034",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00000000",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000002",
  3140 => x"00003574",
  3141 => x"00002c89",
  3142 => x"00000002",
  3143 => x"00003592",
  3144 => x"00002c89",
  3145 => x"00000002",
  3146 => x"000035b0",
  3147 => x"00002c89",
  3148 => x"00000002",
  3149 => x"000035ce",
  3150 => x"00002c89",
  3151 => x"00000002",
  3152 => x"000035ec",
  3153 => x"00002c89",
  3154 => x"00000002",
  3155 => x"0000360a",
  3156 => x"00002c89",
  3157 => x"00000002",
  3158 => x"00003628",
  3159 => x"00002c89",
  3160 => x"00000002",
  3161 => x"00003646",
  3162 => x"00002c89",
  3163 => x"00000002",
  3164 => x"00003664",
  3165 => x"00002c89",
  3166 => x"00000002",
  3167 => x"00003682",
  3168 => x"00002c89",
  3169 => x"00000002",
  3170 => x"000036a0",
  3171 => x"00002c89",
  3172 => x"00000002",
  3173 => x"000036be",
  3174 => x"00002c89",
  3175 => x"00000002",
  3176 => x"000036dc",
  3177 => x"00002c89",
  3178 => x"00000004",
  3179 => x"00003028",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00002e4a",
  3184 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

