-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity VIC20_CARTRIDGE3 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_CARTRIDGE3 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "5104132041EC3184494576544765451D4596441D1675D745916478B80201B113";
    attribute INIT_01 of inst : label is "3441D0450501167441D351449460772521000000364082A0CC81B7B286923124";
    attribute INIT_02 of inst : label is "1930C2096477540535FB722071C71F7A40B716534496DD19E1B02030A82C064A";
    attribute INIT_03 of inst : label is "4A305634308A5585560D05D95113078CDC10E1271D8DE58E40D6ED1841558565";
    attribute INIT_04 of inst : label is "CC94F6964DCB687862A225129761303B964CBDB44850B5645356444D51CB5851";
    attribute INIT_05 of inst : label is "1191D110CA62188E1564E015915626349C12104147B94D1E508E2388E2386744";
    attribute INIT_06 of inst : label is "1DC1551DC5551DC1551D846851D3495535404364D910958A11DA6AB0B0CD1345";
    attribute INIT_07 of inst : label is "4D12449A9B152536015D132D1259CADF48C900CB584075407055477206DEC955";
    attribute INIT_08 of inst : label is "274504D2647654459049761D12868585244DD2121D02C105DAA8905DEE8D0510";
    attribute INIT_09 of inst : label is "1611B6A0D5CB184A4CB184A4346584A58662C0618510D1E589524504D2476544";
    attribute INIT_0A of inst : label is "168904241585555444220158C910400245CD19928AA110478063294880D12244";
    attribute INIT_0B of inst : label is "59011B1065341A0E04C492213082223840888A1D5045A3415535645C91460D5D";
    attribute INIT_0C of inst : label is "C91601113040444D9344407A404500013252E113101C1054501D906184776041";
    attribute INIT_0D of inst : label is "D4A85492A500724706640110493494441916011106040444D890DE06E520D506";
    attribute INIT_0E of inst : label is "EE931044049E12013D1E7759E20BDE751AA1810DA8054D3400704C10D0110168";
    attribute INIT_0F of inst : label is "213445B20583068B958CE13454D5DD0E9DC8479B5725A8B21B764D3470CDC954";
    attribute INIT_10 of inst : label is "747469D59045033001571220410109315C5AA874C5C1B1544854B540106605D2";
    attribute INIT_11 of inst : label is "339874088A28107141807864A21E6B15411475700156122AB05106D7324D9B38";
    attribute INIT_12 of inst : label is "77444D141413514915D950161D0652C52088841788843790194B148943676D16";
    attribute INIT_13 of inst : label is "B34618040D60814B0710E04C49A2C10D90A3174D1D3844E5D1D200451A943474";
    attribute INIT_14 of inst : label is "2A500040168E4A854D2A500624505B01CE0BA898C112511D0458491860101444";
    attribute INIT_15 of inst : label is "1911966740825194446D52410C2AB47291E510114D1C9816A18010168E4A854D";
    attribute INIT_16 of inst : label is "D89855085850D1894E82031C749110E52253B080C491102A9EAA107754844050";
    attribute INIT_17 of inst : label is "2660600152A8B32844DC294DD5144001642A89C0A2465942209265981A850818";
    attribute INIT_18 of inst : label is "55475921350D055544DE15104616256044804616246044904616276044B04616";
    attribute INIT_19 of inst : label is "46186C0499384807975888801FC590104404075D19014B9AE04516BA25150D05";
    attribute INIT_1A of inst : label is "C183B0911AAABAB051A444B46AA9104515144CC11101115110109C4084990788";
    attribute INIT_1B of inst : label is "511D304494451885855811C2188585181801854913044C5111DAA99687746451";
    attribute INIT_1C of inst : label is "25611121CB06322241204A317018D314400544864B44D15245DA15C1119460C9";
    attribute INIT_1D of inst : label is "48A844541F20894EC20214446A8744D15245DA151904834104CD5D5D9DB67477";
    attribute INIT_1E of inst : label is "0864444115159148461624418C4982253B080C511134D1345499768540889C47";
    attribute INIT_1F of inst : label is "89D5115CD541D0120A5D336160119444112B052206A50170210185891631244B";
    attribute INIT_20 of inst : label is "A765DDCD0DDD047746654625442B474429D005A392A1534A9404112D0B08530A";
    attribute INIT_21 of inst : label is "D068834474425645961B44A963898944E43454251846D1D02D18AA01E2A51388";
    attribute INIT_22 of inst : label is "7759C71106AADD90A47472A81414A36D1A46582CAC114145444097619B5408A4";
    attribute INIT_23 of inst : label is "2884418A51622A44044C2745276544AEED10550B796608637DE7512292467D1E";
    attribute INIT_24 of inst : label is "7CC9048C048C3BF37BF37F73BF2E6AEA6159D151D373FB72EA6AE272D98744A1";
    attribute INIT_25 of inst : label is "F78E8000043FC32150079F79E80000C9EFFA000011B7FCB0FE3CDEF3A13F4DDF";
    attribute INIT_26 of inst : label is "13F4C00000E4F43A00001077DC80000D9EFBA000019BE0CA0B5365F47200003C";
    attribute INIT_27 of inst : label is "C6C6C6C6CFFFF6D55F5DFFF400003FFFEE000000000100000000031500600001";
    attribute INIT_28 of inst : label is "3939393939393906C6C6C6C6C6C6C6C6C6C6C6C6C6C6F93BFFFFFFEAAAAA86C6";
    attribute INIT_29 of inst : label is "AAAA8056200000FFFFF0AAAAA0AAAAA055555055555000003939393939393939";
    attribute INIT_2A of inst : label is "03FF03FFF03B00000FF80FFFC0EEA802FFF53A00003FFFDE8000000000FFFFBB";
    attribute INIT_2B of inst : label is "002FF400004BE900000FFE8F55006C00003FF03FFD03B00000FFC0FFFC0EC000";
    attribute INIT_2C of inst : label is "006EBA0000000082824141000087D200001FF400006FF800008FF100001FF200";
    attribute INIT_2D of inst : label is "18D6486359218D58C938918360200A9006D800008401160000666400007FFF00";
    attribute INIT_2E of inst : label is "FFBFFFFFF40FFAD0CDDB76BC75001C8F22F4F00C1890E45401D13F4F40000D92";
    attribute INIT_2F of inst : label is "0000000000000000000000000013A4CE53B90E64F900003FFFC03FFFFFC0003F";
    attribute INIT_30 of inst : label is "0000008080880808000000808080000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000080808";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000200000000200008000000020000000000";
    attribute INIT_33 of inst : label is "0000000220002200000002200000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "5FBA13B91E4B799639ADF177D1F5BAE5A5E6976A66BC5AD5D7469C953FC00022";
    attribute INIT_35 of inst : label is "A78A2BBD42FD556FA4E9D3ECE55DEDF3EAEB439E2A67EDD125EE4CB6FE7DA28B";
    attribute INIT_36 of inst : label is "BFF834037000031FFCE7ED0DC0000EF7838BFF37000030E00E0DFFDE07EFBAF7";
    attribute INIT_37 of inst : label is "C7FC3880827000032AC2E0826DC0000C086381D077000038282EBFF1DC0000C3";
    attribute INIT_38 of inst : label is "0A08AC00003C4C3F6003B00000A20CFF422EC00001420BFEAABB054144108082";
    attribute INIT_39 of inst : label is "8F0484EC00003C843F4203B000005112FF210EC000030503FE40FB82208FC10F";
    attribute INIT_3A of inst : label is "36064D4DA03A4413A4E44849079846FC8A0ED3639100249B15C000010248CF90";
    attribute INIT_3B of inst : label is "22D0271D709D8604B8050C00366199424492D72CF4DE1D13270160C9C0903270";
    attribute INIT_3C of inst : label is "A8000080000EAA80000AAA828202AA800A00004000FFABFF00AA51B1B13900C7";
    attribute INIT_3D of inst : label is "0A95A01555C000258580000000370015A015554AAA800002A20800828A000000";
    attribute INIT_3E of inst : label is "CC95A01555C0002585800000003700153FFF49501415A03609E555A555658580";
    attribute INIT_3F of inst : label is "DCC8D8CC0CC0CC6268B0F2965FCE5E8DCB08E8960047C8C589488115FE9CC5DF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C30C3920CFC4B3CC82784474B66648FE3CF3CA8320F8B2C8F23CB8B28AAB0023";
    attribute INIT_01 of inst : label is "A4A39BD6B76B6F6B5697B74808214A2D4280000CD83D0C10C49BED12CFB07020";
    attribute INIT_02 of inst : label is "764DC430686B6922BB6DB324C30C36F0C8B53855D5FDD252986294A25008CD0D";
    attribute INIT_03 of inst : label is "41C186343D00D20ADD45815555411470905C5225F9CE6C7D48D95528823C01C8";
    attribute INIT_04 of inst : label is "C48ADF38C98B60B6159D0923FED221266584B7DC802E044470444509928B60A2";
    attribute INIT_05 of inst : label is "15929640C999B4015DCF1AA779DC3B389C5909C2DC445613A530421044016849";
    attribute INIT_06 of inst : label is "36420C3E020C3E020C3E04141D234992BA7290A6D924994AB9E9F76254050149";
    attribute INIT_07 of inst : label is "CB22E8FAB6360737B529222D2C164BBEF1C30F8B7080F8A0E0830E926F34820C";
    attribute INIT_08 of inst : label is "3F8F3CB2C4777481294BFED2DD4181C12C8B1BB11A41013F3DD8D3FFDD8D0F23";
    attribute INIT_09 of inst : label is "04710EA0FA4934C184934C083E9B6C134D92883741A9713D0123CF3CB2C77748";
    attribute INIT_0A of inst : label is "110E86204D0158545401125705014A880E41521596A529F6685C05C48A900840";
    attribute INIT_0B of inst : label is "95AF56F3960AB597BA09542693642925A90A49929A5541A592BA569B52C54E12";
    attribute INIT_0C of inst : label is "B60825928298D5A56166A8E58A09AA2B969A9928263498E69A356965956490AF";
    attribute INIT_0D of inst : label is "3AAA456AA9D85D493958A9AA66168A663608259AA8298D5A50A429AE99A429A5";
    attribute INIT_0E of inst : label is "5D8011A0846DDC09BF6FCBF29417FFFF2AA949A9AA97A6B4B410A0246A020110";
    attribute INIT_0F of inst : label is "D11AA98242A20A6766B0101448DADE4D918B49414A25488229B7AD1497454AD0";
    attribute INIT_10 of inst : label is "B64A6559696958C22B5420A966952803549AA95A8ACA8C9C8B56248020A68959";
    attribute INIT_11 of inst : label is "8D667416662498D26FCAE15A529598C9CD9D64822B5420AA92759EE8C0816A00";
    attribute INIT_12 of inst : label is "878489249E6B818DE11622B5028082024010BAAE50AA9E63020809099094AD95";
    attribute INIT_13 of inst : label is "83965A092750C0080A157BA0959E0282508C08452A000C1959D9C0061A9A0694";
    attribute INIT_14 of inst : label is "AA9D34201103AAA456AA9B4BD492982A89B6642F0A551225AC942E596824AC0A";
    attribute INIT_15 of inst : label is "AD168444816B5ED596A69A02401A9A62D2C108100D04DA06A18D001103AAA456";
    attribute INIT_16 of inst : label is "606461A06468958B64C5A830F8E5AD9722D9016A0CE5ADAA19AAA9765A94A4A8";
    attribute INIT_17 of inst : label is "0B7168056AA88C040AD5C5CD968648A3B42AA19EBF4A118155D3A1101AA6A8AC";
    attribute INIT_18 of inst : label is "C30E812DCD3F80C30FB0DD2008190871416008190871414008190B7141500819";
    attribute INIT_19 of inst : label is "09EBA8AE8E64891654B925003ACDA42B590A83CFD6420F03C80C30F12DED3780";
    attribute INIT_1A of inst : label is "45A252A70AAAA6B212BC56AD6AA691490A180849D6A21295EAED56AD80268A68";
    attribute INIT_1B of inst : label is "DD2DC29665A90006465C50450006465C5A0255A92C0430959D9AA9A6A74A4850";
    attribute INIT_1C of inst : label is "21425290480A60016698AFC1BB0D121C48AD9835644A9D6A6D9AE98250A7748D";
    attribute INIT_1D of inst : label is "A6AAA4A8ACF38B6405A83996AA944A9D6A6D9AE9D59A5770D00DDE5E52B654A6";
    attribute INIT_1E of inst : label is "245B65A9595D2A6408190942484DCE2D9016A0A75A9A12A75A9B66BA516C5095";
    attribute INIT_1F of inst : label is "3D6DAD2C694DDC128A9DC041B752A7435298093406A6A0B3900206425921343A";
    attribute INIT_20 of inst : label is "98A116CEC1120784487869084A2B468015E34440EAA915AAA743529A2604FC27";
    attribute INIT_21 of inst : label is "2B6A82C484B28461EBAD8AA840407040100588BA2E8B62EAB624AABBDAA10053";
    attribute INIT_22 of inst : label is "CBF2CFF245AAD562CCBA22AA100423772DCB4854D82108484468E9BA6D9B508A";
    attribute INIT_23 of inst : label is "2ACCA58B3244C149295C3F8F2F774A6D0124A18B5B8215437FFFF24EA9597F6F";
    attribute INIT_24 of inst : label is "BFC333337777AAAEEEE219559D519D1D95555995D040840C40CC08B3FACE80A0";
    attribute INIT_25 of inst : label is "7D1D0000083DE38000014FF0D0000006DFF023F8CEFBCC0EDF330FD300000027";
    attribute INIT_26 of inst : label is "00001D8F83C0000C0000367D0F00000E6DF7C000030BBEF07DE78015181780D1";
    attribute INIT_27 of inst : label is "489DE2374D7DF3FF393CFFF3AA00AFFD4E000010000000000000020000200001";
    attribute INIT_28 of inst : label is "EA95403FEA954000156A956ABFEABFC03FC01540156ABE83FFFFFFFFFFFFE237";
    attribute INIT_29 of inst : label is "FFFFEA02F02A0000000000000000000000000000000000002A95403FEA95403F";
    attribute INIT_2A of inst : label is "07FF033FD03000001FFC0CFFC0C3FF033FF030FF80CFFC0C000006A8023FF530";
    attribute INIT_2B of inst : label is "008FF100001FF200001FFFDC00000000007FFFB00000000001FFE8C550040000";
    attribute INIT_2C of inst : label is "007FFF00006EBA2FF400004BE9000082824141000087D200001FF400006FF800";
    attribute INIT_2D of inst : label is "004004010010042110B10C1306124C2460C008022401B0000000000000666400";
    attribute INIT_2E of inst : label is "FFFFFFC0000F00034578E0A21D03848DA970C4416009C0000000000000000001";
    attribute INIT_2F of inst : label is "000000000000000000000000002940D03EBFE56A40000017FFC0BFC00000003F";
    attribute INIT_30 of inst : label is "8000091919019191800009191908080800000080808808080000008080800000";
    attribute INIT_31 of inst : label is "8000000020000800000002000000000000000000000000000000000000019191";
    attribute INIT_32 of inst : label is "000000000000000000000000000555570000055575455D554000075555400000";
    attribute INIT_33 of inst : label is "C0000555DD455DD5400005DD5540000880000002200008800000022000000000";
    attribute INIT_34 of inst : label is "88AA66A0891A29A06844A8658986A9808068486511998948AA106A969A85555D";
    attribute INIT_35 of inst : label is "9261AA242694251522248A811048829AA886192A4A18A8A890862A64904A0596";
    attribute INIT_36 of inst : label is "7FF400004000010EFFD0D00D0000047FF35FB43400001BDE0D2FFCD29289286A";
    attribute INIT_37 of inst : label is "4FFC7400004202091FF0D20209000004AB0B6209B400001C218DC741D0380343";
    attribute INIT_38 of inst : label is "00000208827F04302822000001F130CD800C00000688333D08B0054144100A0B";
    attribute INIT_39 of inst : label is "0C00000000007C21301213000001F210CD080C000005444B3C84305082DFAAAC";
    attribute INIT_3A of inst : label is "0E8852CFBA034AD3E456487044C504C08D03E444E50008171C400004C002DF04";
    attribute INIT_3B of inst : label is "1C708D3C72D0006434040D4198F127C57F03260C892E11007B00F81EC03E07B0";
    attribute INIT_3C of inst : label is "018AAAC0000401000000300C30CC000030C000A000000155555554055A95080A";
    attribute INIT_3D of inst : label is "ACD62595D92A003CF3C000000033001625973540600EAACC30CC20CC30C00009";
    attribute INIT_3E of inst : label is "80D62595D92A003CF3C00000003300163FFF018C2316259859335CF3557CF3EA";
    attribute INIT_3F of inst : label is "13B2F7135F2F3DF61B50B2231085122921B6FD3BBFE7FF9712602BD901A03114";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "43443B446B2D9146890911008000094E59850B54263985098250B279CAA80C88";
    attribute INIT_01 of inst : label is "A191A77B699DEE0A3B8DEA08BEE80B452200000C94B2E29A2D1DFFB447B69B44";
    attribute INIT_02 of inst : label is "42A26B88380B0B42D1EC9A4451451EFAAD37F24FD3B6828E093452B41621EA98";
    attribute INIT_03 of inst : label is "A90508DA82EE421066525044468A6A432F25E193343CDECD37F2EC29F25A6509";
    attribute INIT_04 of inst : label is "6D0B649AA0D34892400020295DCC8DAA80AD15568AC0929285A92A2802D348A4";
    attribute INIT_05 of inst : label is "A0020A8A200090AECEE4CAA3B8EDF1F207EA1A30EFB8330EEACAB8AE2B8B0B0A";
    attribute INIT_06 of inst : label is "8E52698A92698672698A5743602A200270850409A0230213702DC89426168CA0";
    attribute INIT_07 of inst : label is "1024090001CB5B5AC0202B4D2246D19ECA6AACD348A40894849A63B477FE1269";
    attribute INIT_08 of inst : label is "40904104110000A42690EE022254527640906F3642147643F203243F20329024";
    attribute INIT_09 of inst : label is "8370DE0906D11448AD11448A4090409040A4D07760E730EDA42410410410000A";
    attribute INIT_0A of inst : label is "021A4B4BE48E081818858DA43286AAD04B2026020800276A8680E26D2893220C";
    attribute INIT_0B of inst : label is "8A5F09270849F23BB9162BA24DABA0D89AE83642659185964271A0A882583628";
    attribute INIT_0C of inst : label is "4A8862864464C09AAAA094EAA436005F2A648864D935645965382C800800861D";
    attribute INIT_0D of inst : label is "ED0283380A82800870AA4826AAA909A13A88E282D8464C09A1E12A7E86CD26DA";
    attribute INIT_0E of inst : label is "68048423610A29A091645916AB891451A80270280080922AA85891A1C21A2021";
    attribute INIT_0F of inst : label is "08C0BA9818B8E2A1A243A8580A02C21C88D348092B4D2D0C28909A80A4121025";
    attribute INIT_10 of inst : label is "920A82482C9A0B34A27532881F0B4253E2A2002B705892A6D27CA29E9622E84A";
    attribute INIT_11 of inst : label is "91AA1A42224784C61F37F80A84A4892A6850A2B4A275328025607EEA05282988";
    attribute INIT_12 of inst : label is "8381A8A159FBA6202082D9FE1A068A6ABAAE997EAE997E241A29AAE99C3084AC";
    attribute INIT_13 of inst : label is "9B8800685FE29129A87BBB9162926A30E290C2A42A8A3388686A0A10B81B9190";
    attribute INIT_14 of inst : label is "80A8A862021ED0283380A22A00B458DFE09110A810A8002274B84E2001A17C68";
    attribute INIT_15 of inst : label is "8342B3B0B40A7B5EC0A2A81032E00AB45265365321361BB20C2A32021ED02833";
    attribute INIT_16 of inst : label is "4F4F4EC381498ED262902114F0702AA9B498B40844702880E880AF821930BB09";
    attribute INIT_17 of inst : label is "50C42E206602B0F0492CFA608672D0225CA00EA2B06ACE142010ECEBB826EB4B";
    attribute INIT_18 of inst : label is "1A638A409C63D61A6232002868E051C40C9868E051C40C8868E050C40C9868E0";
    attribute INIT_19 of inst : label is "D2C8817DDCA2D0DC80800022BFA021A4085AD51602126398ED61A63A409C67D6";
    attribute INIT_1A of inst : label is "69BAB41D3200203A02CC09CC0002A948E050F6685253928525FA5CE821024EA2";
    attribute INIT_1B of inst : label is "CC280617A09A113814B10362113814B10B8B819EC0EF018787C00C30BB0B0A93";
    attribute INIT_1C of inst : label is "412252E169A8350DDFE8BA05281EEDA6D2897CA1FB098E67ACC02AD893B3BB6C";
    attribute INIT_1D of inst : label is "BA02BF0D8A20D262DC2117F0A00B098E67ACC02A857F820C26160E0202280083";
    attribute INIT_1E of inst : label is "BA4960BA582E26B868E052CBB67E83498B70845FC289C26399EB300AB40D74C0";
    attribute INIT_1F of inst : label is "0C6C2C232A5E82C41028069E249AB3B052E9A8F9EE06EE2CE12A3814BED9FB09";
    attribute INIT_20 of inst : label is "A882021C1202908008382848084380A300EA8087B40A0CE02A3052EAB86680F2";
    attribute INIT_21 of inst : label is "2A0024108086009255556A008D0838A30781B695A5795C2215C30033E802842C";
    attribute INIT_22 of inst : label is "5916551AB080A02A470AD800ADA89590A4393A21614A760AA29E5695A56AAEA9";
    attribute INIT_23 of inst : label is "625302D15A2B3808C2A6409040000808202182D37F2E800D91451AB2A4009164";
    attribute INIT_24 of inst : label is "7FC37F7F7F7F7B3B3B3F7BB3733BFBB3FB3B3B3F73FB3FB3FB33BFE51254A108";
    attribute INIT_25 of inst : label is "500420B5325F47000000CF78C30FE30DEF30DF7CC13F4C09EFF000000000001B";
    attribute INIT_26 of inst : label is "0000019EFB0000009BE0C000000000024F43000000077DC03FC30000009F79C1";
    attribute INIT_27 of inst : label is "349E38D24BFFF0FF360CFFF0FFC0CFFC0C000010000100001000000000000000";
    attribute INIT_28 of inst : label is "555555400000003FFFFFEAAAAA95556A8015554000000001555555555555678D";
    attribute INIT_29 of inst : label is "55557FA8603FE40000000000000000000000000000006C003FFFFFEAAAAAAA95";
    attribute INIT_2A of inst : label is "07FFFB40000400001FFE8D550053FF037FD034FFC0DFFC0D000007FF037FF034";
    attribute INIT_2B of inst : label is "001FF400006FF8FF80DFFC0D000012A8027FF5340000400001FFFDD000010000";
    attribute INIT_2C of inst : label is "00666400007FFF8FF100001FF200002FF400004BE9000082824141000087D200";
    attribute INIT_2D of inst : label is "00200000800002040118000088442E4304E184938918386EBA00000000000000";
    attribute INIT_2E of inst : label is "FFFFFFC0002FAABEBAA07ADA80C0444FDFF0E88A2008A0000080000200000800";
    attribute INIT_2F of inst : label is "00000080808808080000008080AA952A80154015400000007FEBFFC00000003F";
    attribute INIT_30 of inst : label is "0000000000000000000000000001919180000919190191918000091919080808";
    attribute INIT_31 of inst : label is "C000055575455D55400007555540000080000000200008000000020000000000";
    attribute INIT_32 of inst : label is "0000000220002200000002200000000000000000000000000000000000055555";
    attribute INIT_33 of inst : label is "0000000000000000000000000005557740000555DD457755400005DD55400022";
    attribute INIT_34 of inst : label is "00000000000000000000000000000000000000000000000000000003F0000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "FF38000080E00E0DFFE000020000083BFF834038000021FFCE7ED0E000000000";
    attribute INIT_37 of inst : label is "81D078000084282E7FF1E000022808287FC3880828000026AC2E4826E2F7838B";
    attribute INIT_38 of inst : label is "000011420B7EAAB40000482209FC10D0A089000007C4C37600345054154E0863";
    attribute INIT_39 of inst : label is "2D00001305037E40F40000400001F084D0484D000007C843742034A20CDF422D";
    attribute INIT_3A of inst : label is "FC35152F30C0300C03A83A00600421068C34045500EA8344800000045108DF21";
    attribute INIT_3B of inst : label is "25306B16BBC4215242FF914D01884224084E50920150854D406FC3501BF0D406";
    attribute INIT_3C of inst : label is "024000C0000020C00000300C30CC000030FBFF0BFF100000000000FFFFFF48CF";
    attribute INIT_3D of inst : label is "A8E91A6AE62B003CF3C000000033AAA91A6B3A8006040046024C30CEBAC00006";
    attribute INIT_3E of inst : label is "80E91A6AE62B003CF3C000000033AAA9FFFFE44190691A75157154F1557CF3EA";
    attribute INIT_3F of inst : label is "ADFF144626FC17B2009A0792C35E3D8207CFEF81C0A7F7104040F78354467BE0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "A20A2F38AA2FC208899999A8AAAAAA208A2889E2A8BA289A2E88B8BB5667F188";
    attribute INIT_01 of inst : label is "C84220AD0886A888AA2A8888A0B18B322200000C2096C292CCC689B30A22A3F0";
    attribute INIT_02 of inst : label is "2A968B09B9888B230AAA8B308E28698A0CDA226B9AE222226CB222F2222F33C3";
    attribute INIT_03 of inst : label is "994CE8C9B6C22233230A380002A0CAD3236F311A663F9A973063222FF48A889A";
    attribute INIT_04 of inst : label is "CCCC38AA0ACD8A8B26AA2AA42888CCCCA89FC2088994989889C9CA82A2CD8A82";
    attribute INIT_05 of inst : label is "2AAAA6A2C666C89328A92FCA2288FCFDAF23222F88C8A22B8AD2B0AC2B08888A";
    attribute INIT_06 of inst : label is "2E348A2E308A2E788A2E77736A249661358AC8D426226626260899CDE8324292";
    attribute INIT_07 of inst : label is "A228BA254CC9C9CA56222736A262CCE88A8829CD8A9880488E228BB31AA6008A";
    attribute INIT_08 of inst : label is "88A28A288888889210A2BA2023333A3288A232222233328AE23328AE233262A8";
    attribute INIT_09 of inst : label is "8A228A2622FE28889FE2888988A288A288B3C8A2225222B89228A28A28888889";
    attribute INIT_0A of inst : label is "23210B338C888898988C80AD324C99C886221220002222999984CE0F3F622C88";
    attribute INIT_0B of inst : label is "21022B7CC8C063E284022B210C9B24C846C932201099C846213488A922F3232F";
    attribute INIT_0C of inst : label is "DB04022100208842B088408ACB02FCC6CA122210082720841022304208888AC2";
    attribute INIT_0D of inst : label is "B4548A2952259488CCACB210AB0400882B0402230402088423E3021A2323030A";
    attribute INIT_0E of inst : label is "22C8CCF2B33269124E6398E62B08E38E295233525548404948894322F5222232";
    attribute INIT_0F of inst : label is "488CC2923790AD898A9364CA8922223366CD8888AB362F43A8184248A9323363";
    attribute INIT_10 of inst : label is "988C922230422A7CFD9062AC8A8B2CC4622E009C6B6795A0CD98988CCCDA4229";
    attribute INIT_11 of inst : label is "84CC9BCCCF33308CC2318888C923395A063098BCFD9022808CC22A3949D62A08";
    attribute INIT_12 of inst : label is "9BA8962330A809D22A6A806226C98A46B0AC8418AC8418A526291AC84CC81622";
    attribute INIT_13 of inst : label is "904420C8C622322908CE2840228642332294ED922B09307222694923695C4888";
    attribute INIT_14 of inst : label is "95224892232B4548A295249A6AB228C626C888A92323A98A1888B1108323188B";
    attribute INIT_15 of inst : label is "7A628088BCFEAEAB88A02838332000B3A22A22A22A22A90A029222232B4548A2";
    attribute INIT_16 of inst : label is "73737316767762CD92F3F46134A222283364BCFD10A22280228030998489C6B6";
    attribute INIT_17 of inst : label is "9E8CE4225209B40C94698A066101F3F1A8A012A5B68A023722A2A02369671373";
    attribute INIT_18 of inst : label is "E28B8B36B8ECF8E28AE26624889C9E8CC8C8889C9E8CC8C8889C9E8CC8C8889C";
    attribute INIT_19 of inst : label is "E33863188889CCC9A88000043FD6230988C2F8E2623889A2EF8E289B36B8ECF8";
    attribute INIT_1A of inst : label is "2690B2C22E00008B21888488800024889C9CA02261026222102269A2533008A9";
    attribute INIT_1B of inst : label is "222A4AC88842222727633223222727633908894284DA13222620020889888962";
    attribute INIT_1C of inst : label is "3A2A2222290888DD0A29CB49ED222820F3F6089988946110A000023362808A02";
    attribute INIT_1D of inst : label is "8A01CEBE7A65CD92F3F40088A008946110A0000264288A986C3226626048A8AB";
    attribute INIT_1E of inst : label is "098988C222311088889C9D88A03297364BCFD102228E251844280000B0F34188";
    attribute INIT_1F of inst : label is "122222230232A689252A4D89E16280A1222908C8DA5709E5222227276280CA1A";
    attribute INIT_20 of inst : label is "84166A3F46A248A989B9A8C9889498907A6488CAD15228A548A1222B08DDA40E";
    attribute INIT_21 of inst : label is "04955888AA8AD94608208A558C89B9937358A04220882005C2035562295641ED";
    attribute INIT_22 of inst : label is "98E638E207952A270801915529088C822088AC7322723C84884D09826098AC84";
    attribute INIT_23 of inst : label is "E10816CC222B4AA88CA888A2888888B22AA2B6CDA22B1D8C8E38E2B611858E63";
    attribute INIT_24 of inst : label is "BCC22EEAA6622EEAA6622622222EEEEEAAEAA66222666222EEEAAA7C2A0A93F4";
    attribute INIT_25 of inst : label is "000007DE70015301780C17D1C0EDF330FD3027BFC0000006DFF00000023F8CEF";
    attribute INIT_26 of inst : label is "0000026DF70000000BBEC0000018F830000000000067D0C03DE30000004FF0C0";
    attribute INIT_27 of inst : label is "950FEA540FFFF1EAAF1EAAA1FFC0DFF40D0000000000000001780C0000023F8C";
    attribute INIT_28 of inst : label is "00000000000000000000000000000000000000000000155400000000000003FA";
    attribute INIT_29 of inst : label is "00002AAA45400000000000000000000000000000000001000000000000000000";
    attribute INIT_2A of inst : label is "23FF5300000000000FFFDC000003FFFB000000FFE8C55004000003FF033FD030";
    attribute INIT_2B of inst : label is "824141000087D2FFC0CFFC0C000003FF033FF03000000FF80CFFC0C000002A80";
    attribute INIT_2C of inst : label is "000000000066641FF400006FF800008FF100001FF200002FF400004BE9000082";
    attribute INIT_2D of inst : label is "80C08FE30000002401B00000010044000002110B10C1307FFF00006EBA000000";
    attribute INIT_2E of inst : label is "FFFFFF40001FAAAAAAA48D351E300065555656454881C20C2308308C20C23017";
    attribute INIT_2F of inst : label is "8000091919019191800009191900000000000000003FFFC03FFFFFC0003FF83F";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000019191";
    attribute INIT_31 of inst : label is "00000000000000000000000000055555C000055575455D554000075555400000";
    attribute INIT_32 of inst : label is "C0000555DD455DD5400005DD5540000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "000000000000000000000000000000000000000000000000000000000005555D";
    attribute INIT_34 of inst : label is "00000000000000000000000000000000000000000000000000000002A6C00000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "B43000000BDE0C2FFCC0000003803037FF000000000000EFFC0D00C000000000";
    attribute INIT_37 of inst : label is "2209B0000004218C0741C0000000A0B2FFC7000000202081FF0C2020807FF31F";
    attribute INIT_38 of inst : label is "00000288333D08B0000005082CFAAAC00000208823F04302822000000001AB0B";
    attribute INIT_39 of inst : label is "0C000001444B3C843000000C140CF903C00000000003C213012130F130CD800C";
    attribute INIT_3A of inst : label is "0030000030D4350D43543000000000000C30000000C0030000000000F082CD04";
    attribute INIT_3B of inst : label is "3FE0FF3FF1C000000000000C00200080020C00000000000C000003000000C000";
    attribute INIT_3C of inst : label is "54000000000ABAC000055541050155455540000000000000000000FFFFFFCCCF";
    attribute INIT_3D of inst : label is "0EEA503AAAC000186A400000002AAAEA503AAA85554000005405554400400000";
    attribute INIT_3E of inst : label is "34EA503AAAC000186A400000002AAAEA3FFF0000002A50155545550555586A40";
    attribute INIT_3F of inst : label is "0AF2D3A9A88E1F57A0FF2C916FEE788440451CE2207865BE148ED008F35CBA54";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
