-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity VIC20_BASIC_ROM is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_BASIC_ROM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FCC8FD1C1F989D60DED00019E76699B2BB3E5640626120703410EC35D0DD9B3C";
    attribute INIT_01 of inst : label is "87C919999C705ECCD6A469FDB3699B3C4165049C494406B8912EF76C3BDEB245";
    attribute INIT_02 of inst : label is "393521927FC1F0A9FC6ADE49BC6B26E7133A40CEB09361DF393DC78CD0BC98C9";
    attribute INIT_03 of inst : label is "5181070E460490E2760387642783846930E11A4C46D18653C3C140D82423F462";
    attribute INIT_04 of inst : label is "5B54B07F29B44950741442C1E7F0707291849EE070701A658764074156118E7D";
    attribute INIT_05 of inst : label is "107CF045B91046EC3C398CC5D4443640741E618B7645A435181BE7062544C392";
    attribute INIT_06 of inst : label is "99169090BA447DFCEEC9898AA98BAAABB998746465461C666B4E60E49592F0E7";
    attribute INIT_07 of inst : label is "49889B8650190601913B2649C08749D921400292C6571D97559894554020D6A4";
    attribute INIT_08 of inst : label is "C078C96308E316800F3490D2CD1C37D9E6AC084D48002053988B4188D0002229";
    attribute INIT_09 of inst : label is "7654085C9226E4064EC918C17486764554D3546577502CC51CD148AE08CCA438";
    attribute INIT_0A of inst : label is "0AC28339108515C2136A41D90A432404943243407240351321615C6507041320";
    attribute INIT_0B of inst : label is "6053A8074C1C84714D850921D741340509210A8C044101450D4C891C1023721C";
    attribute INIT_0C of inst : label is "0A6121436143437C41A244564DD34140CD2D20341430354334B50B49DE562102";
    attribute INIT_0D of inst : label is "DDD89F35054408005D2D2C03371147614421C323404B1C4D08374677406440A8";
    attribute INIT_0E of inst : label is "99D9614B045241D2418F142B64E14114F209120902C4B4CCCDCE0041ED2D0350";
    attribute INIT_0F of inst : label is "0414B350438D0CC3A2649916433098C90850A324014526031832144E106CC9CD";
    attribute INIT_10 of inst : label is "824C3010850DC953322B001331403616140AC90134214405D00B04C4DC225430";
    attribute INIT_11 of inst : label is "6418D24914303182C5B89D434465762C2D033A431645451CE0010514924DF34C";
    attribute INIT_12 of inst : label is "41657771888205C33C0191414E340304C5116CD451184C900424B7840388A3A2";
    attribute INIT_13 of inst : label is "80911A89121012680C83015451070C8010860526C98531431A07458956446AA8";
    attribute INIT_14 of inst : label is "144511442C4105A0350441081071450212344CC1186360C027C5C2328C812484";
    attribute INIT_15 of inst : label is "130085D0D0C037C94CF14353A11CF3431484623707090DC413480538B0538D28";
    attribute INIT_16 of inst : label is "DE0C985E104C24DC2143430114D5345073709314F24202A0C8F28322245A045F";
    attribute INIT_17 of inst : label is "D234C63362103489F13747478D2CD9324E2C37873AC1E0CE306518673AC1E0C0";
    attribute INIT_18 of inst : label is "1041C91076727434684444332B4D335013A1501004CA0E0DC98530394418643C";
    attribute INIT_19 of inst : label is "073801CDCD033183440C843049364091A218124413243437274C1C1189304638";
    attribute INIT_1A of inst : label is "1296E355966515771521130321655B84064128CA4E214CC00124C7A31B11BB46";
    attribute INIT_1B of inst : label is "C2014C04269D931737019C31515565CDC50451B3C5202AE8A3290CC401840C41";
    attribute INIT_1C of inst : label is "D991413491498C53070C20524D0453034A900A70516C05094007172BA2A9B22C";
    attribute INIT_1D of inst : label is "041158A3CC1C3174D1355CC0C1E0C1072725243625B633881CDC31C330C51E05";
    attribute INIT_1E of inst : label is "8C1130130D20484120320048423004000C046161904C17474054446010CE3324";
    attribute INIT_1F of inst : label is "301D5DD17300C5009F579093820E081161C918A030C8B84103C808C20170B830";
    attribute INIT_20 of inst : label is "403626868EC91032B20C9D60505242A1072968651123016676710D37744D1D57";
    attribute INIT_21 of inst : label is "35634034A94014C1128C86559101C505D818730CB1C43298B0C704521080100A";
    attribute INIT_22 of inst : label is "34D341D935403441C1044D32614343500370C4C4C1853352405351404DD04D24";
    attribute INIT_23 of inst : label is "556445466091460524005244C8311505525460C105C0004110356D034409374D";
    attribute INIT_24 of inst : label is "5AA3649355A000428CD0D43078CA2B074B4D236614D044091E1E1D914B320441";
    attribute INIT_25 of inst : label is "8D5060951DD207449D8D51929B0444A185020C185450E896C36341250001ED03";
    attribute INIT_26 of inst : label is "14C6C1486329808A80945741D83415346D04AA2645698E65821B08164124CD88";
    attribute INIT_27 of inst : label is "9093745324811B14C00934D04B26C50C11A38D0CE180AC1C000B258A445D18A3";
    attribute INIT_28 of inst : label is "01090A0341C050909090909034930C134918341D92649370080D0524B6634914";
    attribute INIT_29 of inst : label is "40D34E280E401082756454C648A80384324068425D1049C10D0D332434BA85CA";
    attribute INIT_2A of inst : label is "A68C5C861DD61C513403A697771C49E9252DA58C01E1E034588D20A143714120";
    attribute INIT_2B of inst : label is "A264D5DE9E91E0C0818C881929324091271C8104EE89958240B0559046424A43";
    attribute INIT_2C of inst : label is "0D0408A0360A106810CE413404D1CB01158915A9113C612DD119D9521549D03B";
    attribute INIT_2D of inst : label is "20240114B4037643400CA0A37433303009290902CC94170A8550016420CA0D2D";
    attribute INIT_2E of inst : label is "38200154120140B1151760482B34E248511778D1342203A26402841108210074";
    attribute INIT_2F of inst : label is "15527893C60CA86100C10404184EE192AA1B28CCE04602418320E0900E018ACE";
    attribute INIT_30 of inst : label is "014815A8B0C8014217667660331405910AD30426F010BCE141010F0114504133";
    attribute INIT_31 of inst : label is "925440441889B8ABA2801CC95176491D3544119D1211331061314001A0076212";
    attribute INIT_32 of inst : label is "E2A3A0A1A08745754747776766764262EA86855DC522B898958999DDD1115551";
    attribute INIT_33 of inst : label is "2544D58320C39000314C438AC83F1EBC010022EA66686010600502132030018C";
    attribute INIT_34 of inst : label is "AA667774445554406733CA264D9064590547646CB320456031040450107C4D31";
    attribute INIT_35 of inst : label is "0000C6338A2408060C04D9274CC510040531455924676664D9064590C922098B";
    attribute INIT_36 of inst : label is "A81F0999DDD1115552222B89A05085121100023302214A1AC5504C8838E38A14";
    attribute INIT_37 of inst : label is "99025499D927491254328C8600E0805924664D9064590C93154477664C2F01AA";
    attribute INIT_38 of inst : label is "8D11244512244204104A22458546D92D193058DA51508730B14248468C092116";
    attribute INIT_39 of inst : label is "5CC9280147648D55186240C01501099A19005215A50764812144D890511D3044";
    attribute INIT_3A of inst : label is "061810A1A30C04D4AA312A84895273394906000C2C0D09858DC3016270C4D0E0";
    attribute INIT_3B of inst : label is "4801C318449356205387040BA5A58C50E9FA72D091240A4A6100526486D99000";
    attribute INIT_3C of inst : label is "DF747115D4520434188D2532269926D8D49158C101A886A220C4D88310576045";
    attribute INIT_3D of inst : label is "4599D9C90E91555690422B449010D48000876C43498637613003674288802799";
    attribute INIT_3E of inst : label is "1438C502AAAAAAAAAAAAAAB001F203F3C2FFF803F300F2413203A00041444D04";
    attribute INIT_3F of inst : label is "24CC11833401092D6872067BFE8A077849D98588D20096038C30C09032700A13";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "57476757B2020FA1C330EFE4A0219769BB80001BABA88B98B9D0B99F48203052";
    attribute INIT_01 of inst : label is "06C56615413D87CD34C541353446D375744E54E14E116735D172CF5E3B8AA8AA";
    attribute INIT_02 of inst : label is "4DE534C783097DC00C44101ED3F373EE147F660376057553CD321C312DF1E01E";
    attribute INIT_03 of inst : label is "DE45171F7914E1F74407C4957747C79D31F1E74C791E4B33D356D66157480314";
    attribute INIT_04 of inst : label is "63DC7177D1799C4317E111C5C4D179931521E0D179919C4DC495317E731E4782";
    attribute INIT_05 of inst : label is "9CF0F4373444797F3D1E12132C49449317EC620F8998005E5120041077510557";
    attribute INIT_06 of inst : label is "BE44B0E0304CEF0133031122230302232110300001334F985F935155D5E7C170";
    attribute INIT_07 of inst : label is "4E80A6622288498919A424690A8661D98458222A40E50390E4389020EAA0842C";
    attribute INIT_08 of inst : label is "C0AC06C029B02984A93A0092412F04711EA0C001445AA21914896A2014853061";
    attribute INIT_09 of inst : label is "667680D0602518902101960B76877B5776CB544747011096284D849C08099403";
    attribute INIT_0A of inst : label is "491EB5D0220F38C030442210086A024C008476534188B0EA77444F3D54898276";
    attribute INIT_0B of inst : label is "A0EA6422A89C0E71AD0A4A90A2A864090E83AA6901CE424A4ECD429424B3903D";
    attribute INIT_0C of inst : label is "A58B044777546574C2734B74A98A22C24CACA3325882316B30743649E93B0343";
    attribute INIT_0D of inst : label is "DED4293A4BC9C0545CACA4B03341579156928032B084288A4427B67A6074AAA2";
    attribute INIT_0E of inst : label is "11E5E3CF1A9A629A6A422AABA4224124900E920EA2C9BACD0E41D741DCAC8302";
    attribute INIT_0F of inst : label is "3A3A9080B1F7002E426698A62AC280080DD48266C8A9A78E3801288823B3114A";
    attribute INIT_10 of inst : label is "41B0B02899D999D5C361176C00AB6667772999C8300460D29A3F1808AED2A70E";
    attribute INIT_11 of inst : label is "66A49A69A6BB5C3C8E889EC24864B714D949266A16566A287E022EA69A6920A7";
    attribute INIT_12 of inst : label is "52855791540B3A801F914293A71F8C088A107C64A23C80292622556641438242";
    attribute INIT_13 of inst : label is "BCB0460B05443194CC9A32168503380A30AF2DB7C29922301415555554554619";
    attribute INIT_14 of inst : label is "20280A00181102607445440AD55357235705244540FF8B0003B515E20C486CA4";
    attribute INIT_15 of inst : label is "270A42ECAAC23A4A419380430320A2053CCDF3293A2602042208E106F391C9E4";
    attribute INIT_16 of inst : label is "21099DDB3397841EE647531004E23BEC806B903A9032825140A23012A49928A6";
    attribute INIT_17 of inst : label is "9106B900703AE442D30683F8483CAF20810F06C207CE7001F083200207CE7000";
    attribute INIT_18 of inst : label is "7202999B96909714A6810D026689005303030304089951D9999921444BA114E8";
    attribute INIT_19 of inst : label is "672FCE418009C05473C088A068B62C8B02A4DFCC2267654666F0E4220DC33A10";
    attribute INIT_1A of inst : label is "228A7E4390E4393D0BAF02092654BA0095A6A9784226480043410F1353353D80";
    attribute INIT_1B of inst : label is "9B0BC40A861E7C351A337B034374A2024288D2C082A9099095D3000D9BCD000E";
    attribute INIT_1C of inst : label is "D5DB6DA69A61A9F0182C0E1861965E28611A0D7BEF70828288093626426B7124";
    attribute INIT_1D of inst : label is "3BAEBCE37061C183E5B94C880A4D480A67082A2B38B80E0CACEEC00CC00D22C1";
    attribute INIT_1E of inst : label is "2D12213340E92903347F84D41B744884CD04935555481495A09496EE91780C20";
    attribute INIT_1F of inst : label is "2C9955953243CFC45E97AAC37AA72A596BCF3CE0300AA355FF44480041457CFC";
    attribute INIT_20 of inst : label is "CFF806A00CC0CCB152AC5E14281ADD63744454DD20EE02A67B4300E565699953";
    attribute INIT_21 of inst : label is "314350747744030A19408A55D201060DE4640200A00403743B00085D2004200B";
    attribute INIT_22 of inst : label is "B2CB22C5B1407699226606A64447475110BB08C886553092A86A90B206DACC96";
    attribute INIT_23 of inst : label is "350D60E0EA5960259682DB77B8E01A08717CF00154C000998075A9256012B72C";
    attribute INIT_24 of inst : label is "4683168315041810B4C49113417CC1072B6C931516C081411D1DDEDB6D243888";
    attribute INIT_25 of inst : label is "CC596A1129C837061C0D1A50662241121160209A9C9C9111332B22A2A8D28CAA";
    attribute INIT_26 of inst : label is "340D0A6A6A0452AA8034A729C1169996610A6816054189151A58C88465C74CA4";
    attribute INIT_27 of inst : label is "C2DB40FF74012F19FA29A65A6F0B4F0812E040178D02982C2DC0474056119450";
    attribute INIT_28 of inst : label is "50455403ABC0F0CACACACAC8269BB0236DB89699CA729A6498A4A63297036DBC";
    attribute INIT_29 of inst : label is "051BAD16A5D855404444457840560754A09046011D86020945CCB04476540111";
    attribute INIT_2A of inst : label is "457014199129907135044774591445110A1D11DD051950B4944D029554605006";
    attribute INIT_2B of inst : label is "4046151DD111D0D44181C450A0A0200900148949110116802082990A64282800";
    attribute INIT_2C of inst : label is "AC0ED86075C60458517444B006DBCC2595BCA66C994C99519219DC5A654DD004";
    attribute INIT_2D of inst : label is "6E80270A900149617241194046A07142A0A0A00981155F05055A8902A211ACAC";
    attribute INIT_2E of inst : label is "D020A9461AA96AD314179002AA1073C4A21797E0906DC84046A981172AA04810";
    attribute INIT_2F of inst : label is "08715FF14E0991140B0212901609151A4446667040B50523800B0E00840B4100";
    attribute INIT_30 of inst : label is "106CA6146F0B328AC775796C9F088994094008096040980D65A40525945555E1";
    attribute INIT_31 of inst : label is "514490A85455454460682401108442510954615EA020136011928410140B9744";
    attribute INIT_32 of inst : label is "C04051617047857957947847857941551101C12E418045544A71911915D55D51";
    attribute INIT_33 of inst : label is "184AE12C03890000451142A1246829F0002CA5111110141A9228644445445517";
    attribute INIT_34 of inst : label is "5565565676676688A8C2FB0681A1685A066554A4AC2C86F29208082823AC8A92";
    attribute INIT_35 of inst : label is "C0044193400A0BCBE7A4E5176B0124EC41B24190A4B7574290B42D0411128665";
    attribute INIT_36 of inst : label is "AC2BE919919D5DD5D8312677722409A2975176064064B2064118B84B2383422B";
    attribute INIT_37 of inst : label is "5D040601E580605815047899404F01108494210942504119D6564545574BE1AA";
    attribute INIT_38 of inst : label is "014A04900415129015458D44554AE18121E020E9606B0B1060418A4538062194";
    attribute INIT_39 of inst : label is "EC8B60095446355128954780212601112589A1282B27A852A073E058541EA152";
    attribute INIT_3A of inst : label is "2EFC2A83436DC058D81236C80DDB4377BD8B0700144A8A8ECA4001B3A004A454";
    attribute INIT_3B of inst : label is "8002DC04A153B81482FF388046678022BF6FFFB3D2A02B6ABC05A2B6B1D5DF2F";
    attribute INIT_3C of inst : label is "1D857A55EA50013A248EB8402DD28AE4A8AB438A336CCD83038C20CE32B5A8CE";
    attribute INIT_3D of inst : label is "88282A8AAC8260BAD8A336A0E828E14C448BA513AE4D3BA856ABAB9280C48761";
    attribute INIT_3E of inst : label is "2420C2F2AAAAAAAAAAAAAABC0BF300F202FFF80FF802F1033183A00002088E81";
    attribute INIT_3F of inst : label is "170021A3380020177A8EDE4F635791AA05E5418AF280EA2AC58380EF33640CAC";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "7646466748BAA6697570547038BA01111367A9A60231012312043231030400AB";
    attribute INIT_01 of inst : label is "50101044440104114115114045101441001015095010504005857C825F5DB5DB";
    attribute INIT_02 of inst : label is "50004404141400155111541007F401AA45400614060504040045404141010590";
    attribute INIT_03 of inst : label is "0025549000950904116420100424200049080012004024081020240640901019";
    attribute INIT_04 of inst : label is "5402094404451058000108250509411854511509411941012010800000802014";
    attribute INIT_05 of inst : label is "4102060440420000818054104215410800011920110452200544458040116200";
    attribute INIT_06 of inst : label is "0901020845200002100221032113321033213321032100411010488011040980";
    attribute INIT_07 of inst : label is "FE2D1115F4571434A6D0D2B6B6A9A866F302966430484100C0312900EAB80100";
    attribute INIT_08 of inst : label is "D8862E48CE18A8ED80B8B208642CA0B82E009A3C11CABE9B9AD1C489C19CA6B8";
    attribute INIT_09 of inst : label is "0929308E1B4AAD26D81A623A9BAA3AA22971A2A2A1C846038A20E1CEF8ECC282";
    attribute INIT_0A of inst : label is "2E08031B5A04C222962242A92A936C27B2622A80386D14F0A23B8C3198E40529";
    attribute INIT_0B of inst : label is "F470BB6347070C15B0103EFCF34B8343C7C383002C5C1C961CB2780F8DBF0430";
    attribute INIT_0C of inst : label is "A461B3322AB33BBA920A0AA09A9262D977270C54610D5581DE10AAACEC3743D1";
    attribute INIT_0D of inst : label is "0C2180B8A920B36147270628DC0913851A84A3860CE18A9831B3AB3A9930847A";
    attribute INIT_0E of inst : label is "8ACA0823A8E382E394238A988108A42D0BC73F470CE0BB327C508CD8472795DC";
    attribute INIT_0F of inst : label is "0C0E1E14BC828E0B8739CF33C005F21F2CC383B8A08208E6823860E69B808822";
    attribute INIT_10 of inst : label is "2841B622CCEECCE307994C2048AB33BB30EEEED4FA8003A2AC83A8ED001F0830";
    attribute INIT_11 of inst : label is "3942CB2CB28031A230420EDB0AB09946AA387BB4DB9BB08A20A38238E38E3884";
    attribute INIT_12 of inst : label is "9D2182BD10AAE0A38886140C058820CEF0868EA30386BD82C2FC0088080AEB87";
    attribute INIT_13 of inst : label is "921BB9A1B220B41A142948681A27965946A18208EE0048C3985099911A91A8A1";
    attribute INIT_14 of inst : label is "85C1705C96442A7B2199EB222A8E28462872C15CB2729010AF4AAA59A5039A23";
    attribute INIT_15 of inst : label is "83EC52CF2DFBB0221608958B812538A4967219F3E0D8783F38A229903A8D6302";
    attribute INIT_16 of inst : label is "86ACCEE1888C6360330B878DDAE8BA6A8D882B400AFC8A692D388384A1206585";
    attribute INIT_17 of inst : label is "0858C0A594230E32F8D8E329A28EE386242C982990EA5A560880222990EA58E5";
    attribute INIT_18 of inst : label is "4812EE06838E00C0B216D23B30E085BC4B80A85A4ECC2200EE0048010A62220E";
    attribute INIT_19 of inst : label is "53842E163322058884528E380F33CBF0960210EB3B308803B80383382278419A";
    attribute INIT_1A of inst : label is "39982307C1F07C0DC3F5896688A03DA2A08244C2308012321051604807004021";
    attribute INIT_1B of inst : label is "28A02B06A88E704B4BE48C38240020705ECE0208E2022CC1E31BE332E4628ED8";
    attribute INIT_1C of inst : label is "888A28A28A242008E2EE28A28A28A5862A8A0E80208E0303530541B307A015E5";
    attribute INIT_1D of inst : label is "AAAA863881C70614CAB29ED65861204BB861E1E1E24031A2A1C205670CE020AA";
    attribute INIT_1E of inst : label is "90A415A4650ACAC84A61AA42C102505651B0AC88A212AAA884A8AB3298C23074";
    attribute INIT_1F of inst : label is "9E00A00A780AE0064ED3BA3840A580A2A823863A48E818AA73E1416A0A223642";
    attribute INIT_20 of inst : label is "E738DA223EB9B14E842E8EA123AE886AAA221A0026258AA2B29C650082A020A7";
    attribute INIT_21 of inst : label is "54AE07922A90941A4C0E800002565850E18F5B4E8561380080358E0038AD3968";
    attribute INIT_22 of inst : label is "14514252148B2066391012513BA13ABD050010B0142299860AAD84169264F508";
    attribute INIT_23 of inst : label is "1A0680C0FA082782084820094D59A8528E8218EAA9E006440698828001A25945";
    attribute INIT_24 of inst : label is "B005480548B08259895225B498C29969C9971D484072FE1C84EA0E082381E0E0";
    attribute INIT_25 of inst : label is "158A28CC20724968E526EDB713543EE2CC09C16247650ACC494142A261222500";
    attribute INIT_26 of inst : label is "CA947A9A847B2E980891A1C8788A0641858A0048122C10CAA6A1237383101501";
    attribute INIT_27 of inst : label is "38209A00016403A9038E382083B8E0924239A68C69A6EB2FB41A200BBAEEDA68";
    attribute INIT_28 of inst : label is "7912A9CBA9620A1212121218B2C803382082082C330CE3962D0301CC80C82082";
    attribute INIT_29 of inst : label is "3EEF0092A4032208686868C61A64BA9E440FB21ECA6138D0303B3A232002A888";
    attribute INIT_2A of inst : label is "2101C1E664244F78E07A22A90BD234882684EE002CCEE5809AF26AB333070570";
    attribute INIT_2B of inst : label is "862964600AA84561587E51CB2B2ECDB3EFD2F416AA18A20AC71646B11AC2CACA";
    attribute INIT_2C of inst : label is "0B23126BA926999E78C61B6CB288208A298119A1618E44EE42A4634826F028AA";
    attribute INIT_2D of inst : label is "42A4A7881A89090505288B8739078716AB2B0B21688AA0AE1CE6D76C0E88AB2B";
    attribute INIT_2E of inst : label is "128211924AA92A3AEB633DC900DA58E383A390C75A41268629A9A6678067155A";
    attribute INIT_2F of inst : label is "D29E9439E0ACCEE929E3A52CA21CA8A72B33B9C148CADA78239062B234A809A6";
    attribute INIT_30 of inst : label is "6EB3AA939C14B5662A223292619AF2072078CE206A521A6124A727861A44AA59";
    attribute INIT_31 of inst : label is "6A20A60B23A2A2A28694923830E0C3830E0C3C6CE8EA969E1E8F3086908B22A1";
    attribute INIT_32 of inst : label is "2A86868687B33A32A32A32A32A32AEAAAA3A182C3AF6AAAB09C8AA8AA8AA8AAC";
    attribute INIT_33 of inst : label is "9A08EA404DADF000F33CCBB17C85317000992333333117E8AEC8684C4C4F0E8C";
    attribute INIT_34 of inst : label is "AA2AA2AA2AA2A958040505A96A5A96A5BA22209E40526A7A69AA26259B926669";
    attribute INIT_35 of inst : label is "2022BA7A0BC979271CA3CAA29C1825971A5EAA8B202A222C8B22C8B288947AAA";
    attribute INIT_36 of inst : label is "012418AA8AA8AA8AAA4EEAAA0E2DF986228628629628BBE9E8AC96F4946A09B9";
    attribute INIT_37 of inst : label is "8AB2689ACA2689A268A216223269AC8B2022C8B22C8B288522A2A2A28C642C00";
    attribute INIT_38 of inst : label is "58B1602E68E2CE2CA2285232220ACA28286A23EA8E9CD6B73EACD26C96B349B2";
    attribute INIT_39 of inst : label is "81D148AA222140A8A822B16B8AA1E8882AA8587284A3A1AACE9CC1ABABCE062C";
    attribute INIT_3A of inst : label is "841EEE69858723AD468F59E1746D859906C8694EA13838383853B42E14E18381";
    attribute INIT_3B of inst : label is "3322406B8C83686A884592DA23B962E2A7A9DF5C4EFC919071EA84198A88A7A4";
    attribute INIT_3C of inst : label is "85EA17A85DA22C34E30D2B94C442CAE303258964959E94684D66E5759B939A6E";
    attribute INIT_3D of inst : label is "48101EF2BA01206A6C86DA838FC0FE9C388B02C34A1437A380028B047353A17A";
    attribute INIT_3E of inst : label is "6BDA664AAAAAAAAAAAAAAABC0BF40BF0007FF007F80DF803F141300222048D30";
    attribute INIT_3F of inst : label is "91A16E69B8005F0BF16E472ADF777CBB28CA3A1269A22685E245622486962270";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "CCCFEEDDCCEDDFFEDED0DFCDDFECEDEDEDCEDDDCDCCFECCDEECEEEFCDC5555DD";
    attribute INIT_01 of inst : label is "5D5D75575757577575D55D57555DD7575D5D755955D5D5D75C7DE7DF75C71D75";
    attribute INIT_02 of inst : label is "5D7575D75D75D75D75D75D75D6ADD7AAD5D7565776575D755D5D75D757575595";
    attribute INIT_03 of inst : label is "75455515D515515D55454555D545455D5151575455D54551536565565595D759";
    attribute INIT_04 of inst : label is "7554515D555D5551555D514575515551557557515551575545551555D5154555";
    attribute INIT_05 of inst : label is "D5545455575455D5151557555455D551555D5145555D544557555515D5554455";
    attribute INIT_06 of inst : label is "01550050554014ECCCCFFFFEEEEDDDDDCCCCFFFFFEEED5D55D5551155D555115";
    attribute INIT_07 of inst : label is "211FDDD9BE662726361C98C63B9DA27608B07E1230D8C360982363B0BFE85540";
    attribute INIT_08 of inst : label is "E2B0E6F0F2C39B4C7D1122D3C22F0B22CA20492332367367B0CD9892332348E2";
    attribute INIT_09 of inst : label is "8588B0B0D3F33FC883210F28D89CB488847989888989B02D34F7422EF8466D01";
    attribute INIT_0A of inst : label is "2607DC4B9F08CF027888B122286FCB23220888B9C34C98E888888E388B86C989";
    attribute INIT_0B of inst : label is "B3ACDBF3BF3F08ADC237330CE3BD80EFFB02FDA22623233A331073233FCFC022";
    attribute INIT_0C of inst : label is "922C0888888888BC32E08488422CA2F4E6A68C9E238C9CBCD9988896E73A02BE";
    attribute INIT_0D of inst : label is "2D233D118BC6233336E6FCC1D8888B8C096F412ECC4C34FB325B49B4848899B9";
    attribute INIT_0E of inst : label is "6446E38F29249165630F096863E382AFD23AF33ACFE69CC0FFC075B666E68D8F";
    attribute INIT_0F of inst : label is "C9CA08CACF9F0405C99626C9BD4C62762223CD9B06965B0C3810EC4E3AB522EA";
    attribute INIT_10 of inst : label is "D35338212222662C4C88F5D4BA94888888F26630BC59A223239F284F7C7CF915";
    attribute INIT_11 of inst : label is "94B065924971C4823BB86EF58D98D8B0222C99488C8C8C34E7811A492596F0B9";
    attribute INIT_12 of inst : label is "B8C888F88897CF413D4DEECEDE3DE484BC0DBCA3B138FF3FCFD88888888825C9";
    attribute INIT_13 of inst : label is "B0C19FCC19988CF87F67D59B662E3004F81E124BCA66E3510C88480084884000";
    attribute INIT_14 of inst : label is "59B66D98BC6626D1999B462D5988D8C8D88DA32362D4F5220BD666E3CF3DBCB3";
    attribute INIT_15 of inst : label is "0BC031DE32F0774200D08C8B822FC30E3CC0E1CCCDCB7B73130E4C08F08F8E78";
    attribute INIT_16 of inst : label is "3E16622C38B1232C48988F80C9CC08208CB1F3CFD0AFCAE38FC3910FE238873E";
    attribute INIT_17 of inst : label is "D0CBDC3C8C2F7830E0CBC38B8C3C2E0CD22F0BCC0BC2E132C182222C0BC2E043";
    attribute INIT_18 of inst : label is "E3216620888CC8C89B1000119BCD0C90CB82C040C46666666666E19888A66D70";
    attribute INIT_19 of inst : label is "5471EE32362C4099B5FB84F1B6C9B76C8EF0C7C3119999999B533313C2F39F3C";
    attribute INIT_1A of inst : label is "1286E58260882208C32D0BCD19982B8248512B123E19B8323055455154055545";
    attribute INIT_1B of inst : label is "670786ED842DC4C5858DB91199D443232B0462E3C26427736C4B9200038C04F3";
    attribute INIT_1C of inst : label is "65659659659256E0DCDE056596596C189326E9B1E5B07A7AE6EFD89DCD885DE0";
    attribute INIT_1D of inst : label is "8820B8F392BF4EF9D6B5B8323BF78C8598CFEDEFCEC6178EA3FC4B0F48422056";
    attribute INIT_1E of inst : label is "AE0DCDCB0E69B98801D7426269B83F372C188C9999B85F9E8BD8D8F54B1214DC";
    attribute INIT_1F of inst : label is "3C216216E088EE446B9AE9F3D69E1965A78F38F0AC493966C78373758999BCD6";
    attribute INIT_20 of inst : label is "CC78C0B22EF762018FFE6E62237266E19999B8722D6D0999118B8E4405A1016E";
    attribute INIT_21 of inst : label is "DD8CCCD98888BD330184A2642AF23332E33EC3848B021088B12C0462109F138B";
    attribute INIT_22 of inst : label is "DB6DB266D9888B66E19B2119889988BDCDF137FF3766788CD5B1C9FFE16277D8";
    attribute INIT_23 of inst : label is "26099090A9659E165989240B97D3A8AD81B8E0459B802966C9944259B26119B6";
    attribute INIT_24 of inst : label is "9BC19BC19898B0E3DF722E3C8B120B95B946CDD8DF623333662224249F0BCC4C";
    attribute INIT_25 of inst : label is "2765A766226DC99F262721FDDFDA367222C1F25A665F3266D1ADB161110226FC";
    attribute INIT_26 of inst : label is "C9F7A86860912A28889889A2625A65996D08BC1B0626F3652A5B4311BC7527B3";
    attribute INIT_27 of inst : label is "F165BCE59B828F2B5F1659659F2BCE382AF38F3120AF2F2F0D699888CA3230E0";
    attribute INIT_28 of inst : label is "F19998CB97C2E16D6D6D6D6499671311967859666D9965BC6C96DADB99899678";
    attribute INIT_29 of inst : label is "2213514BF229998898989B12332E19B48CCD9B26659833F33336F99998889666";
    attribute INIT_2A of inst : label is "8B13333666266FE0CCCC88898BFC33222266226622222F4AB08225888888CC8E";
    attribute INIT_2B of inst : label is "C88466666226627327233232E2CCB02C0BFCB73723221108BCB0652D94B0B888";
    attribute INIT_2C of inst : label is "D62E7CE19B8E19B4D312251899678E165B16D9E66DB866226166566906F46488";
    attribute INIT_2D of inst : label is "F5589D09B8488C8CCCD224C8844CCCCC62E2D223C2266E132211F88A4E2266E6";
    attribute INIT_2E of inst : label is "78626599665599F29A9F69C86DF4E3C3311BB1D734F788C88467866D19A629F4";
    attribute INIT_2F of inst : label is "ADA1B9F3CE16666227C10A488B26221189999BD3E056F6E38135E6223E188B8E";
    attribute INIT_30 of inst : label is "8DCF9999BD3E0B8D5995B5B8D789F45226F0C426F122BCE492622F12492266E2";
    attribute INIT_31 of inst : label is "5598BCC5999999999D88B4263098C263098C265D18DD913816B3D88D98875998";
    attribute INIT_32 of inst : label is "25CDCDCDCDDB59B59B59B59B59B595555577261DE73111110716566566566566";
    attribute INIT_33 of inst : label is "B9A976D40F0C480A308C208886489D50024FD11111320268FF049888888988B1";
    attribute INIT_34 of inst : label is "449489489489482A1E4F9D1B46D1B46D188888B8E4F8EED1D3BB4EED3AB0EED3";
    attribute INIT_35 of inst : label is "0009F7D18B843B0D7D50D659BD369000250D96629A19958A6298A622227D9444";
    attribute INIT_36 of inst : label is "0F6D6676676676676B339111082032C81D8DD8DD8DD8BADF8670B07E31E18BBB";
    attribute INIT_37 of inst : label is "66589A244689A2689888B066326196629A18A6298A62222F58989898B12E4600";
    attribute INIT_38 of inst : label is "372CDE08DF14BEC88895F5999988D6A626C122E18DB1FD393D96FD98B05BF662";
    attribute INIT_39 of inst : label is "32CD8899999BD266A2599B82B65B86458696E03DAD1BA04B1DB1D2637276CDCB";
    attribute INIT_3A of inst : label is "1C7431F1C11E506F7F0FDFC03671B5175708118453333B333B210DCCD8433363";
    attribute INIT_3B of inst : label is "23B2C4D8B66388108B1F3429988BCE605B16C8B163148140D41188DB56656C1C";
    attribute INIT_3C of inst : label is "6C59B166C46A263B238EC980E6630AD230118B8D3DFCF7F00F4EA03D3A9BB0EA";
    attribute INIT_3D of inst : label is "882821E3C282608A7080D8B33F38E6B333A36663B237392D9BFC474AC0C2DB16";
    attribute INIT_3E of inst : label is "D9F8E2C2AAAAAAAAAAAAAAA00BF005FD08FFF00BFC0FFA0EFA80300922088E30";
    attribute INIT_3F of inst : label is "1B0256C3A80204BF515421BC4914440896D63625F3026F1BC28F426F01BC26F4";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
