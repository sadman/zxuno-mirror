-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity VIC20_CARTRIDGE is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_CARTRIDGE is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "77721DB6C6F16AAC8DC8A9318844A088891E951D1551913389195191C241B1E1";
    attribute INIT_01 of inst : label is "0391788C02905506406451A5044114D03414141B74040610E4E9393934E38D22";
    attribute INIT_02 of inst : label is "100A004766744819040D19267645103841D03801110354D4240E13540E03744D";
    attribute INIT_03 of inst : label is "40434642262AC2476491DD1044346475744E1C901181522B8344410344028419";
    attribute INIT_04 of inst : label is "85A6C9411091204424614244A05891D5104634434581559E2654657072404605";
    attribute INIT_05 of inst : label is "C9C1DE1545E12470617168A35D954519D02D10D1344114D23665368D9120DA22";
    attribute INIT_06 of inst : label is "774435C2B4E275DF72144491DD181D18199816D19494D037D344C346768DF441";
    attribute INIT_07 of inst : label is "650770441515C9C1DE10441725451051347CD1A2476640650D05DD34899DDCD2";
    attribute INIT_08 of inst : label is "53427600470440002BFE851E24DD35220491D01D10199016D5981D011344CC35";
    attribute INIT_09 of inst : label is "3578995D524644D41D81D0C00778CC102019D5E24576658464D5111D5340111D";
    attribute INIT_0A of inst : label is "1456145601D81D95011D38DD99D251D46571C530DD990000003D000F25789959";
    attribute INIT_0B of inst : label is "81DC1D05D81D0474D113778D18D8D41D1174D10D05515A544E24626047741456";
    attribute INIT_0C of inst : label is "6891D991376627788260740450074044AA49963B91758EE01D054244AA49981D";
    attribute INIT_0D of inst : label is "4678995D91238D92244DD909DC20981D011810D12475441191DDDDE2891D9E36";
    attribute INIT_0E of inst : label is "9D19C057371554448058D5D912449D12147174090CE246564524656458541B35";
    attribute INIT_0F of inst : label is "99C01103F275DE70D199A30C14405352670441064D9248C3048B46254C559591";
    attribute INIT_10 of inst : label is "244099D4D1CDCD92111999134672488C6247781DDE0766448259409D104104D1";
    attribute INIT_11 of inst : label is "5240660642488CE933824777492802407607675789257674802407607404884E";
    attribute INIT_12 of inst : label is "952742516414B456524003FFC9575D7354A148990198196149599E2656665248";
    attribute INIT_13 of inst : label is "D53126495266305351649CDE237845D89D051C92466549099066491995262641";
    attribute INIT_14 of inst : label is "7495D9A334789D599DC3665067074EEC912CD195D9265D841D90D9E0D5349149";
    attribute INIT_15 of inst : label is "9410000155BF36C14D818DC5112036653664A04D994D9EE38A24066076427627";
    attribute INIT_16 of inst : label is "410D09C9C552449504104108100CD81D053778044150670074246347899C2640";
    attribute INIT_17 of inst : label is "276470A04E04D30C2A8D007441441462744174D0446666055414911251545516";
    attribute INIT_18 of inst : label is "5767144A4495090DD148D99515D32654506714507714038599D1E36478199D1E";
    attribute INIT_19 of inst : label is "5911A24416034780541D50D685D095CDCD1419D9C1145D3C51D9958289D77972";
    attribute INIT_1A of inst : label is "2091918150D1A4824666064278141349100423360724469D99951845289E156D";
    attribute INIT_1B of inst : label is "C119D811011D05C19901D8D020451766724504346075B820D5D5992549244113";
    attribute INIT_1C of inst : label is "6066492346625B21DDE077786484665876467065707670724514C119D811D105";
    attribute INIT_1D of inst : label is "3C83044881849258001000092C009D0992464902A051E289E77936D199412110";
    attribute INIT_1E of inst : label is "1251D320912438900DF679A507464630C38E746449C538C24330902F70E6CEC2";
    attribute INIT_1F of inst : label is "8E38738E210C38E4B46454E2C626C57AA0012C04046382D90E91B31474130CDC";
    attribute INIT_20 of inst : label is "0DE01DE02644104109A255D74A112346448B0E0930189D19169CCC08690D3898";
    attribute INIT_21 of inst : label is "7501094E247774667891DDD191E247774667891D9D191B1491E17447644581DB";
    attribute INIT_22 of inst : label is "459104019A0445CE1491D16419211524091111A705006584B8475194732A4B30";
    attribute INIT_23 of inst : label is "1D1E247464747891D191D1E24746474440089CA4506060202107707507707434";
    attribute INIT_24 of inst : label is "74144462865A2864A284492501904883410E11593449D1541537499147891D19";
    attribute INIT_25 of inst : label is "408008554418199198A6194DD59C20021551060664562AA38667107822055A08";
    attribute INIT_26 of inst : label is "9A3474EAEAEAD190441D934D1114D5411DD1774516740000000000253E43A43A";
    attribute INIT_27 of inst : label is "8D08F08D082449F30D137CD134D1D91268D28F28D28F28D28376545474F565AA";
    attribute INIT_28 of inst : label is "6064562AA386771078222C07707D5959800081515D017382204405CE088D08F0";
    attribute INIT_29 of inst : label is "FEAAAD055FC001CDA12FF015AAAABF5480085441819198A6194DD5DC20021510";
    attribute INIT_2A of inst : label is "000000000000000000B9672F7A85709A429E749259CBD916E66DC6DDDDDFFF14";
    attribute INIT_2B of inst : label is "00C4F13408000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "00000C0000003F4300C27F700000000000F5707000E0B1340000000000FFF070";
    attribute INIT_2D of inst : label is "7776000000003B00000000027776000000003B0A0AD80E7000039FC000003DC0";
    attribute INIT_2E of inst : label is "F13498000000370277761D00000000000000000277761D000000000000000002";
    attribute INIT_2F of inst : label is "00000300BFECD0000000000000030011B583000400000000000000FFF07000C4";
    attribute INIT_30 of inst : label is "FFE3000C3C00000000000300FFF4D033D000000003800002758C00000FD00000";
    attribute INIT_31 of inst : label is "F4C0000000978300B3F8D033D70000000380000EFFCC000038F000000003000F";
    attribute INIT_32 of inst : label is "00000011B58000040003002D6380001CFACC000033F700009783000FFEF3000C";
    attribute INIT_33 of inst : label is "FFF40033D034000000000002758800000FD0300000000000BFEC000000340000";
    attribute INIT_34 of inst : label is "D73400000000000EFFC0000038F030000000000FFFE0000C3C03000000000000";
    attribute INIT_35 of inst : label is "E000001CFAC0000033F73000B580000FFEF0000CF4C3000000B58000B3F80033";
    attribute INIT_36 of inst : label is "00000000E028A000248008000D000000000000FFF60000D573FCC3FFF3FC0025";
    attribute INIT_37 of inst : label is "9CFFFFFA5CF0F002F18000E29CFBFCFA5CF05002F182F8E29CF2F8FA5CF3FC00";
    attribute INIT_38 of inst : label is "00000003AAAA8003D1F00000BF8000000000000000000003F0003F02F18000E2";
    attribute INIT_39 of inst : label is "00000002955680C00002C30000000000007000008F8000008000000000020000";
    attribute INIT_3A of inst : label is "0BE24000000000000000000002A24000000000FFF60000D573FF0CFFF3FC0000";
    attribute INIT_3B of inst : label is "20802000000000200FE0400404C01800000000080FE2400000C0180000000000";
    attribute INIT_3C of inst : label is "00FFFF00002200020002C000000000400D60000800000000000000182D60000C";
    attribute INIT_3D of inst : label is "96CB685299EC8595447742D5767866754765467675445470D591D5151D3891FA";
    attribute INIT_3E of inst : label is "554A83581DD1D0B8100138008120B3C91C034230B18B2043895CA7894145E3B2";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "F05AFC056AAFFFFCA1096180614AB74B892C111E12599232C5259992E0CB00D2";
    attribute INIT_01 of inst : label is "20114544201255884804521104620AE1380C0E2BB8080A281BC6F1AC5BC5BC5A";
    attribute INIT_02 of inst : label is "A80D137675A488D2B50D16B775AD10200DD0204DD2324A93340C02740C126481";
    attribute INIT_03 of inst : label is "5151A4C22000407858161602A4384785B683C8D8A5C212365274AD436A0340DD";
    attribute INIT_04 of inst : label is "4D08B64690B6A0A40A5142C84170D5D100851A738475D1D514B5744C23629708";
    attribute INIT_05 of inst : label is "0A42E124A2100A5272714B306E19A29D5225285A95658A5634B4150592245422";
    attribute INIT_06 of inst : label is "5766373D4730421392249CDE5D902D58AD9098D9D82C64142969336755052A99";
    attribute INIT_07 of inst : label is "762A70B4D2DD0A42E110A7370949949934A3D23C785B52B50D8ED2B58DDDD8D3";
    attribute INIT_08 of inst : label is "2A426520B60A555555554D23C5E15B24DCDE9C2D54AD9C98DDD4A9C2D9A54337";
    attribute INIT_09 of inst : label is "175452D5FF5A40246986208A85844CA2A0DD9D5377654B57D49DD2D92A5BD2D9";
    attribute INIT_0A of inst : label is "25F92579021C219242220FD9D9505F14E941460CD9D955555596AAA5375452DD";
    attribute INIT_0B of inst : label is "421CA1869C62149B123184412C6C1C2221A412424A96E6480A24B27088682539";
    attribute INIT_0C of inst : label is "8C1E1EDA9758094C5352970A531790A4994696E671A5F99C291491A499429821";
    attribute INIT_0D of inst : label is "675452D5D9620D6636A5D6825314D4A5C2905469058780A9161ADA6CF161E835";
    attribute INIT_0E of inst : label is "69927E490A2A648892601211284022920A51A48B20C34B756D34B756DC2057D7";
    attribute INIT_0F of inst : label is "D9509276A05217A0D5D93D84496A7180A5095E96529B58622489C836A0A99A95";
    attribute INIT_10 of inst : label is "0493D1D8EDC20E11D1D15173776048A4816B8416613747489063FC2DA28A28D5";
    attribute INIT_11 of inst : label is "B362A70A5248A8C54580786B6B0FB362B708777545BF77458B362B7085148A80";
    attribute INIT_12 of inst : label is "922490B0A4968A562A7776AA81986EA37832C49DCA902982C9D9D514B6765258";
    attribute INIT_13 of inst : label is "5AC12649224A1090A3A498210384069465C298924A64A9896A64892992A724A9";
    attribute INIT_14 of inst : label is "609D9DA20B5452D9D9337B62A70A49902DD8699D9D0621AADDE0BAB2529692C6";
    attribute INIT_15 of inst : label is "24D55557FFEA3A80A2828E42522436763A66B1CD9D8E9C6CFA362A70A790A53A";
    attribute INIT_16 of inst : label is "828AC28AC2936ADFE8A28A000000E8ED370984348D234B30A60A43A5F527D488";
    attribute INIT_17 of inst : label is "2774803100CAE84A2AAAF2BA43C83C908A51A4B3C899993E5824920191A49625";
    attribute INIT_18 of inst : label is "474628444611C206D858D1D116D20786A2A70B50A4043E89DEDAA177A89DED2A";
    attribute INIT_19 of inst : label is "ED2141A61442CACA4A952A55025825C506982E590298692312D1D1FCF1485ED3";
    attribute INIT_1A of inst : label is "24EAD58210E108929B660A42703CF2CB2000002A1A08459D9D92154A289C525D";
    attribute INIT_1B of inst : label is "4AE9982D02A98D0A9D829CD1236918A67195260B70A62F60BEDED9A4A9A48121";
    attribute INIT_1C of inst : label is "62856163774062216E10598484B74463647A62A440A462B08504CAA9582A9949";
    attribute INIT_1D of inst : label is "F8DC1844CFC8A0604AB24A0CC03295A9FC4B7C12C0F210C1E87E8ADDD1CA1D1B";
    attribute INIT_1E of inst : label is "99522212DAB6800A01CC73A2874B4812100EF6B780002CE04381297C4109DFE2";
    attribute INIT_1F of inst : label is "06D81186022100CC36B680B00F05C71FFDD1210100A8CADE04DE0D148833F0E4";
    attribute INIT_20 of inst : label is "02106212267301A9A93C6A18AA69636B6888400F0C345DAD2C602CC5421F10D0";
    attribute INIT_21 of inst : label is "844324430586B6B58C161ADEDA30585B4B58C1616D2DA700D2B35B597A4BC9E0";
    attribute INIT_22 of inst : label is "ADD6B40ADD85F47304161ED1F521FDD1F5217DB4C132B4FC805F5FD5C32B4030";
    attribute INIT_23 of inst : label is "2D230587B6B48C161ED2D230587B6B48CA0888B6A03030303318728408408835";
    attribute INIT_24 of inst : label is "380484A24D9224C9224C8122A168644AA00812123E8FE0E8360D8361F8F161ED";
    attribute INIT_25 of inst : label is "00A0A815422A055058A528A65504292A05508A81541629514941018CA3084604";
    attribute INIT_26 of inst : label is "D3C6861111111211447DD04FA298E0FB211E3C4830F800000000003FEAA95540";
    attribute INIT_27 of inst : label is "831811831836AD3C4DAB4FDAB41211A84F30C10C30C10C30C15B4484760C4FAA";
    attribute INIT_28 of inst : label is "A8141629514979318CA22883B04313D01800A0505E0694CA28001A5329B31811";
    attribute INIT_29 of inst : label is "C0FC0C0EA555011A8096AA9502A54000A4A81422A05058A528A655E42A2A0508";
    attribute INIT_2A of inst : label is "00001555555540000ACE415CF12889D050134B17505716440787D8872D85DF00";
    attribute INIT_2B of inst : label is "00C3F0FC5088222222888A22220888220888A222222088AAAAAAAAFFFC000000";
    attribute INIT_2C of inst : label is "00002E020080B72700E43F9000EABC0000E6071C00C7F0FC00EABC0000FFF31C";
    attribute INIT_2D of inst : label is "DDCAE80000003B000000000DDDCAE80000003BBFEDD9ACBC0000DF0000003CC0";
    attribute INIT_2E of inst : label is "F0FCA8000000370DDDCAEC00000000000000000DDDCAEC00000000000000000D";
    attribute INIT_2F of inst : label is "00000D22F44EC0000000000000030003FF3B0000000000EABC0000FFF31C00C3";
    attribute INIT_30 of inst : label is "FFFB00043E00000008B60D036FFAC00BC000000000C00027F41E000054000000";
    attribute INIT_31 of inst : label is "F4C0000000E4CD035FFBC0032400000280C000073FEE00000C7E0000B603000C";
    attribute INIT_32 of inst : label is "00000003FF3A000000030031B0C00007FFEF000038E30000E4C3000CFFFB000C";
    attribute INIT_33 of inst : label is "6FFA000BC0B0000000000027F41E000054001C0000000022F44C000000B00000";
    attribute INIT_34 of inst : label is "24B00002800000073FEE00000C7E1C00B600000CFFFA00043E03000008B60003";
    attribute INIT_35 of inst : label is "30000007FFEF000038E31C00C6C0000CFFFA000CF4C3000000C6C0035FFA0003";
    attribute INIT_36 of inst : label is "F2EBF21EB20EB2EAB257B25D70028002000200FD73E000C533FCCF6AA9FC0039";
    attribute INIT_37 of inst : label is "3CFFFDE29CF0F0269CF000EC3CFFFFE29CF000269CF3ACEC3CFFFCE29CF1F4EB";
    attribute INIT_38 of inst : label is "AAA200035555C003E2D00003D1F00003FF80000008008001F800BD269CF000EC";
    attribute INIT_39 of inst : label is "0000002400001860002F49000000000002D00003CDF0000340C0000000C1C003";
    attribute INIT_3A of inst : label is "5FFC000000000000000000005FFC0000000000FD73E000C533FD8F6AA9FC0000";
    attribute INIT_3B of inst : label is "10C00C00000000053F8E800002400600000000056FFC00000040000000000001";
    attribute INIT_3C of inst : label is "FAFFFF0DA41B000B4001180020C00200FB0408049080080001800200FF0CA000";
    attribute INIT_3D of inst : label is "188950A29EC8A606548792D5C783797948447A57A7A4A5B89692DD592C2C52FF";
    attribute INIT_3E of inst : label is "FFCA8330D152CE7030C500820E24108E34D28B1490401062C528A449428E1322";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "5AAAABFFFFFFFFFEACD3AE470B0830D2E922888E420C82FAA020CC82EB2C0CD8";
    attribute INIT_01 of inst : label is "8B8FBB228B8ECC0BA2E3C2CC84F289CABAAEAF2B39C1422C00155AABFFC00155";
    attribute INIT_02 of inst : label is "666AAAA2A1A0A1866BA4E669299AC98AAA898AAA829609AAA26AAAA26AAAA0AE";
    attribute INIT_03 of inst : label is "DF8CAAAB4B8A68183A0E0E8CA972C28393AD2E434710786296219AE9199AAAA4";
    attribute INIT_04 of inst : label is "458AC238E906E72B42BCA40A4CA24747842C4A8F2E856568B091D1FAB90D1C41";
    attribute INIT_05 of inst : label is "F4D4ED8092DA42A6A4ACACC82309E2A479452182D79E497D9092DCA5AB4372B4";
    attribute INIT_06 of inst : label is "08084B33ECD82F0AD480AE42242746B7467BF242490B4B82F482E90909208C20";
    attribute INIT_07 of inst : label is "90D0840A0220F4D4ED9C294940ACE1CE80A402C028391E0A247C024B64242F28";
    attribute INIT_08 of inst : label is "2C9608540AC2B906FFFFE02D02709D492E422346B74677F24247425028AAAE90";
    attribute INIT_09 of inst : label is "81A2C242810AA3C3CA32EA92A4B63E984A060689090B08A80182022024A40220";
    attribute INIT_0A of inst : label is "A33AA3BA76A32A02146EB44A4AB82709EAAA6BBA4A4A1AC6C6FFFFFF81A2C242";
    attribute INIT_0B of inst : label is "F2AB2A7CAB2EB0A4C2AC3BAC210BE3AEBF2AC230308DE80A3A808C8D1AA2A33A";
    attribute INIT_0C of inst : label is "B20E0E42E90A52B6993D2B42ACB3842AAA34AB2A9F2A88814AB08C2A8810A16A";
    attribute INIT_0D of inst : label is "A1A2C24A4ADAA42D90BA4254AEA64B4A90AFE32A8083A32A020E4EA300E0EA90";
    attribute INIT_0E of inst : label is "2AD2B34840C2A1AD0FCA0220E4A102A8CA8F2AD342E909939690993B6307E821";
    attribute INIT_0F of inst : label is "47BAD23FF82F0AE24B47C26BF6CBEE341F527F6D7F7AF69BFED262A4B10A52A9";
    attribute INIT_10 of inst : label is "84B843438310783B1B3173C90D3CED222948B6922D8585AD0CCA03069A69A64B";
    attribute INIT_11 of inst : label is "B90E0C43DEED2A200908083927B0890E1C42595A2C9D1D2F6890E1C42DFAD222";
    attribute INIT_12 of inst : label is "92A4AC0C2EB90AB02EFE97FFE09C23993ACAE3B438350FBAA16D68B090D3FEF6";
    attribute INIT_13 of inst : label is "EA0F60E92A48C42C273E972DA4B67CA34E30AFBB4BC4B37D2EA4AD2F124C74BA";
    attribute INIT_14 of inst : label is "A64646BBC1A2C24646E9190D1841A44106412A464682F0AE64690EA9C27B92B4";
    attribute INIT_15 of inst : label is "036E4EB3FFFFB26892223C30E94E90D0E37D8B243438F2A34990D18413841871";
    attribute INIT_16 of inst : label is "A230303030A90B68269A69A28A23C30692C0B690A42908C4184295AA0C2930A3";
    attribute INIT_17 of inst : label is "A910A2AB2E392BAA8008240AA40A43840A9F29040A888842B9EA028C0C2A82A0";
    attribute INIT_18 of inst : label is "3939C3BB39EC90F8A7B64E4ECE8EB1B0AD1A41B41A7AD26E46429B93A6E46429";
    attribute INIT_19 of inst : label is "E42885384A243AA709EC2FE210E3027E92AB46AAD0ADCAA4C24E4EB300BC2BA9";
    attribute INIT_1A of inst : label is "4102671075CB2924098C43DECA41041028A288F05043AED61692B80B43B202C4";
    attribute INIT_1B of inst : label is "D42A2102742A7254A234A32A4908D099C52DFDC19418A8D90E4E43609AE4A96A";
    attribute INIT_1C of inst : label is "FE05D3D90D0CCA4922DA48B62D048488280A9D2BAD2BA42F3BFA542A2342A272";
    attribute INIT_1D of inst : label is "22C0C19A82ED04CAD2B4212B3ED98E7AA04A8AB49900DB20BC2F884343B8B1B4";
    attribute INIT_1E of inst : label is "AAC8EA40425ABA31208C2382D9190B4AEBA9D1938A2CAA991408410019509889";
    attribute INIT_1F of inst : label is "EA2AAAAAB4AEBA8C9193B2ABEB91200FFA5A4E8584ABE042224EF2F23AFA03C3";
    attribute INIT_20 of inst : label is "A2DA22D8D2A48E1EDAC02709E02AD9090A93AEB3F33124242242012111908606";
    attribute INIT_21 of inst : label is "AB2FABAD82839390B6020E424AD80839291B60E0E4A428B282AA0A1A2A0AE8EF";
    attribute INIT_22 of inst : label is "BA42EA90AA9E6B0DBE060EAD205F5AAC204F9AABAF9C2B893ADD374EDF8AAFA6";
    attribute INIT_23 of inst : label is "E46D83839191B6020E4246D81839291AD2AD3EAB2909290928CA8CA9DA9CBA90";
    attribute INIT_24 of inst : label is "788180B4449B4748B4448A4EE0648D409122020241902419024190640B40A0E4";
    attribute INIT_25 of inst : label is "56A520620EC918838D282890A832A9481883B24620E34A0E8A0CBC3E0A608B48";
    attribute INIT_26 of inst : label is "6C0089202020020A0D266A900EA1C6B0288E5A09A63B1B1B1B1B1B1555555555";
    attribute INIT_27 of inst : label is "6CB6DB6CB69096F3A42DBC425A022024B0CB2DB2CB2DB2CB2A09808819DC3F80";
    attribute INIT_28 of inst : label is "2460E34A0E8A38AC3E0A4D0788370FD80182A1E3CC2FEBE0A844BFAF834CB6DB";
    attribute INIT_29 of inst : label is "C0FC0C2C000000000000000000000002A52060EC91838D282890A8E2A948183B";
    attribute INIT_2A of inst : label is "5555400000003FFFFA80114104FF88110D04004044504441101014F94FA47300";
    attribute INIT_2B of inst : label is "80CFF354660F943E94A50FE943CFA53E90FA43E97E94F5AAAAAA55FFFEAAAA95";
    attribute INIT_2C of inst : label is "00003CC300CB434100C24D8000FFF70000E843E780EFF35400FFF70000D573E7";
    attribute INIT_2D of inst : label is "EEC5DC00000000000000000EEEC5DC0000003B7FDE399EF000007F0000001D00";
    attribute INIT_2E of inst : label is "F35421000000370EEEC5D400000000000000370EEEC5D400000000000000000E";
    attribute INIT_2F of inst : label is "A8002C3BD02F00000000000000030003F0350000000000FFF70000D573E780CF";
    attribute INIT_30 of inst : label is "FFF50000D8C0000034D32C0BFFD700327000000000700031F80F000000000000";
    attribute INIT_31 of inst : label is "790000000CBD2C0B3FDD00014000000318700003AFF7000000D8C00CF8C3000C";
    attribute INIT_32 of inst : label is "00000003F037000000030007C07000039FF50000047900083D03000CFFF50000";
    attribute INIT_33 of inst : label is "FFDF003630C0000000000031F80FC00000000E00A800003BD02F000000C00000";
    attribute INIT_34 of inst : label is "40C0000318000003AFF7C00000C9CE0CF8C0000CFFF70000C9C3000034D3000B";
    attribute INIT_35 of inst : label is "C00000039FF5C00004790E083D00000CFFF70000790300000CBD000B3FDD0001";
    attribute INIT_36 of inst : label is "71D571D571AB712D710D71AEB00FF00FC00740FC33FC00C533E95507879C0007";
    attribute INIT_37 of inst : label is "5CFFFC6C3CF35CEC3CF000E15CFFFF6C3CF000EC3CF0F0E15CFFFE6C3CF000D5";
    attribute INIT_38 of inst : label is "55710000000000FFFFF00003E2F0000003C00000BC00F8007FABF4EC3CF2F8E1";
    attribute INIT_39 of inst : label is "00000090000006180050240000000003FFF00003EEF00001FFFF0003FFFF4003";
    attribute INIT_3A of inst : label is "2FFC0000000000000000000027FC0000000000FC33FC00C533E95507879C0000";
    attribute INIT_3B of inst : label is "0300010000C008001EBC000001000000008000001FFC00000000000000000000";
    attribute INIT_3C of inst : label is "FFFFF5003007E00F0000070200C2400068B400000040010010C209007ABC0000";
    attribute INIT_3D of inst : label is "12D148B4DE2D34B230A3B45CE78839390911392293A0A0BA8E8600402AAA02FF";
    attribute INIT_3E of inst : label is "FFEA8BE24CC2E2BEFB69A28AAAAA9A29AAAA6BA68AA9AEAAA0293761D4FCD8B4";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "55555555555555559EFF5D0B4B89A9CEC622222E2222E292C22222E29207F1D8";
    attribute INIT_01 of inst : label is "B38FB324B38CED23ACE3E8EE48C244DA11999C2840AC9E700000000000155555";
    attribute INIT_02 of inst : label is "52CEA3BBB9B89EE13A02D538B54EEB0A8EEB0A8EE27B84E83AC2A3BAC2A3B89E";
    attribute INIT_03 of inst : label is "8C8C0A073B0A4488A9262A4C08FC8B8A899A6822B23B27FFFFF84E8094B3A8E2";
    attribute INIT_04 of inst : label is "888A523726233BCBADBC9888CCA022224CC8C08FCA926268089898ACA08AC8EC";
    attribute INIT_05 of inst : label is "E7E349084090AD8C8C8CA9A0A629A02227322273084104290A88C89227332273";
    attribute INIT_06 of inst : label is "8888CB16A5A0A629B348A821222233A233A3A2222232BB0A50A2B0888A128A22";
    attribute INIT_07 of inst : label is "88AC8EC92322E7E3490ED8C88C92223248A522A4A8A88ACA0227210A42222F24";
    attribute INIT_08 of inst : label is "3088C8CAC8EDAC53AAAA922A4A629B3968212233A233A3A2222EB2FB280A4B08";
    attribute INIT_09 of inst : label is "49A0226294849373723081FA78243F8189262681898888E93232212210A92322";
    attribute INIT_0A of inst : label is "4AE24AE2302382223B8829222280A228A2B24A2C222238F90EAAAAAA49A02262";
    attribute INIT_0B of inst : label is "38230267230808A5226CC8D2223F230839C92223232B888939088C8EE0A84AE2";
    attribute INIT_0C of inst : label is "A8262A2318AB8DA8A08AD8EDA54B8AD933272B4CC9CAD33E32488AD933272302";
    attribute INIT_0D of inst : label is "99A02266669242A908C62A236B2822B63B632302488A9302222A26869262A90A";
    attribute INIT_0E of inst : label is "12A296888C8C989CCE89212290923024C089C9FFE2E585984658D98C63332959";
    attribute INIT_0F of inst : label is "2AB1A242A4AE2BA42A2AA6C2BEAA8AC8E88EAD2AADAAA4B3E9CE8268C232A12A";
    attribute INIT_10 of inst : label is "78A12E22BE232BEFEDEEDE80B8BF9CE4278C24E30938B89CCF8A52B28208202A";
    attribute INIT_11 of inst : label is "808AE8ED8D9CEC200AA498A8AE69B08AD8ED999A02B9999A4B08AD8ED8C9CE82";
    attribute INIT_12 of inst : label is "62588CCCD9844088319556AA9298A69099A203622BA3B6A24A6668089A998DA4";
    attribute INIT_13 of inst : label is "2B4F8E962588CAFAF9D96F093C242723323B6F658DA8CAE731989616A1289CC6";
    attribute INIT_14 of inst : label is "A06666B28DA0226666B0A88AD8ED977736770266664AE2BA62A62EB3210B62A3";
    attribute INIT_15 of inst : label is "3361BCEAAAAA76C440923F3327380988AC84B202622B22869808AD8ED98AD89D";
    attribute INIT_16 of inst : label is "9233333333248C2960820812492272B25B8C2458962588CAD8AD8C0A12284893";
    attribute INIT_17 of inst : label is "3888AC92494406CB155B78C098898A88C089CA2889777789F8D9224CCCC92248";
    attribute INIT_18 of inst : label is "8888CC8C8422232B10A422222E290A887ADBCDBED8C986C22A22B088AC22A22B";
    attribute INIT_19 of inst : label is "6224C8C8CA88BACC84223323332332F2F02E3172FB6E7265222222B692B8AE80";
    attribute INIT_1A of inst : label is "3231323B23F22CC8C4E8ED8D898A28A2249248BC8C8C9262A262488B33622222";
    attribute INIT_1B of inst : label is "231323B2231332633223332735888C5E8AE8E88D8ED8AD922E262AF84ED89227";
    attribute INIT_1C of inst : label is "8AFB4E90B89F8B3E30938C242FFBBB8B8B84A8CCA8CCA8E8CAC9231322313232";
    attribute INIT_1D of inst : label is "6CA48C8DB60CCF89FA7E262B6493E13EA78A5B23B2289282A8AA822E2E2BFED3";
    attribute INIT_1E of inst : label is "232083CF210A64E62E8BA28308989BCFB24889888A0B2CA00010010010018888";
    attribute INIT_1F of inst : label is "886092083CFB24B88988ACB24800401AA5573B0888A64626222297CC20829373";
    attribute INIT_20 of inst : label is "109130909CA949F1CEA4A629A502908899CEC922862322222240400004101000";
    attribute INIT_21 of inst : label is "0A880E0A0B8A8989A82A2A2A22A098A888AA82A2A222292C22B0A88999AA02E9";
    attribute INIT_22 of inst : label is "C22309E723FACA1A242E2A394C8E72394C8EB28AC93DCA9CE488A62A8FF8993C";
    attribute INIT_23 of inst : label is "622A098A8988A8262A2622A088A88889F89FE88C6636363634C08C08C08E2048";
    attribute INIT_24 of inst : label is "B88888B3888B3A89BF888BFF12109F3C4222222289A2288A2288A2A8AA92A2A2";
    attribute INIT_25 of inst : label is "019CA8840A8A21022FC028412222672A2102A288408BF44C888888E467CC8FCC";
    attribute INIT_26 of inst : label is "2A4A480000002224861114A20C237892A20088A22899C61B6CB1C60000000000";
    attribute INIT_27 of inst : label is "4B24B24B244842A6C230A92109212210A9B28B28B28B28B2848088488488AE95";
    attribute INIT_28 of inst : label is "28808BF44C88B888E4673C8B88A22B88001992022D288A466480A2291A5B24B2";
    attribute INIT_29 of inst : label is "C0FC0C240000000000000000000000019CA880A8A2022FC0284122E2672A202A";
    attribute INIT_2A of inst : label is "555555555555400000010001010010000040010040004000400411555001B700";
    attribute INIT_2B of inst : label is "00D57D0000A5554055555155542555402A555400155505555555550001555555";
    attribute INIT_2C of inst : label is "00003EE700F42F20000396B000FFF1C000D1434D00D57D0000FFF1C000CD334D";
    attribute INIT_2D of inst : label is "BBB92E000000000000000001BBB92E0000003B0505199FC000003F0000000C00";
    attribute INIT_2E of inst : label is "7D00040000003701BBB900000000000000003701BBB900000000000000000001";
    attribute INIT_2F of inst : label is "0FE03001EA44000000000008000300227A400000000000FFF1C000CD334D00D5";
    attribute INIT_30 of inst : label is "FDF000006B40000033FB302CF5C0001E90000000003800007E0C000000000000";
    attribute INIT_31 of inst : label is "0000000034F0300DFFC0000000000033EB38000073D40000006B400CF8C3000F";
    attribute INIT_32 of inst : label is "000000227A43000000030033E0380000FFF800000000000C3C03000FFFD00000";
    attribute INIT_33 of inst : label is "F5CC001AD3400000000000007E0CE000000003000FE00001EA4C000003400008";
    attribute INIT_34 of inst : label is "03400033EB00000073D4E000007A430CF8C0000FFDF300007A43000033FB002C";
    attribute INIT_35 of inst : label is "E0000000FFF8E0000000030C3C00000FFFD300000003000034F0000DFFCC0000";
    attribute INIT_36 of inst : label is "9000160018400400D01450000E014001000000FFF3FCD7FFF3FC000055540033";
    attribute INIT_37 of inst : label is "9CF1F407D241F4E15CF0A0E59CF7FC07D24000E15CF0F0E59CFFFF07D2400000";
    attribute INIT_38 of inst : label is "00000000BF800000000000007F400003FFFFC000F4007C0017FF50E15CF3FCE5";
    attribute INIT_39 of inst : label is "000000C0000003016AA9400000800000000000007F40000000C0000000C00000";
    attribute INIT_3A of inst : label is "41C18000000000000000000000410000000000FFF3FD70FFF3FC000055540000";
    attribute INIT_3B of inst : label is "0400000020C4100205C180000000000000E0240241C180000000000000002000";
    attribute INIT_3C of inst : label is "FFF5000004030003000000000000000000C000000900000040C4000205C08000";
    attribute INIT_3D of inst : label is "E2CC88B3662CE8898899B368998898B8A8889999999A88A426262222282C22FF";
    attribute INIT_3E of inst : label is "AA9FCA61622284E4824B28A2C828B2C828A2882892CA2882C22CCA46E3E790B3";
    attribute INIT_3F of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
