-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GAL_HIT is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GAL_HIT is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "001B11C001B01EE803F15AA8330FBFC2BFF80BEBC1656F9425402A65BFEBFF05";
    attribute INIT_01 of inst : label is "01C049878595512001000B114BEB55523957032A9993A1BDE7DB3C10F57A14ED";
    attribute INIT_02 of inst : label is "14557B766B62000016F5D45126138580D00C9C009BD555C20004D55561AC9700";
    attribute INIT_03 of inst : label is "4445511011100054033C00FFC033C0F3C3157EC000DF4FFCC09B12EAAB0032AB";
    attribute INIT_04 of inst : label is "6A075554200006C9BF60840FE34000E855510E57910012EEE3E0B56155015555";
    attribute INIT_05 of inst : label is "BC3047AF111BF0FEA4ABFE9947E07D05C504550E3B55470000D5F185355116A6";
    attribute INIT_06 of inst : label is "C4CF4000115414004010F6F290440400400CD4140F050C01150C0F1A01054FF7";
    attribute INIT_07 of inst : label is "F80002A8813E59AFE32E2541B3B9010699051A039063C555080D063E8DC01BC0";
    attribute INIT_08 of inst : label is "A38582C000282FCE8C451195A9578687B00077D73B5F8B14B9BFF5B1547D554D";
    attribute INIT_09 of inst : label is "ABF3F8D838955558848A9D0000B1F3E4F3C0EEAAAFC3CFF3F018CC390CCD9554";
    attribute INIT_0A of inst : label is "F4A42A90DA5EBECAB8CA43CF0144CF56B0C03C04F5511AA44283D7E0015436BB";
    attribute INIT_0B of inst : label is "D9011400C8CEE403ECC925AEFA1A00BC50A4B4500A706EAA16CC1024D7C07117";
    attribute INIT_0C of inst : label is "0F93CF03BAAABF0F3FCFC06330E4333655528E160B0000AC70FD01040166A913";
    attribute INIT_0D of inst : label is "CFF3F3FEB0F0C40256A529FFC20001435CFFC83CA79013555535072F70000207";
    attribute INIT_0E of inst : label is "3CF03CAF30480ABEF1A4F75557E20001E355EE4D6E890010015902D403C033FF";
    attribute INIT_0F of inst : label is "ED002DAB8E46ACCA0050400044445101000066BFB942FFEA5B0A84FC0FFF3C30";
    attribute INIT_10 of inst : label is "5536E418D54DB007039C064AC55557A3E9C55200000C336014FEA910980C1C54";
    attribute INIT_11 of inst : label is "156A90FD5B6532800979574D7C463BFBC857780039FA0800023C3FD3D44698D5";
    attribute INIT_12 of inst : label is "D34008B38C05000B55582001581DC55F023E355239A9BAB400B1AA4BED0B45BE";
    attribute INIT_13 of inst : label is "A314BF5F50006A9A5CC15574A959E5BD45AB19384000000B185555D0ABDD00DB";
    attribute INIT_14 of inst : label is "0028EAAD001BE4C9160AA6801A2C0394156F57C0AC53980033C3900B1A3D9B9F";
    attribute INIT_15 of inst : label is "EE2FD66BFF97713E8CDFCE0005CD5557802A78C86F5289130B0905FF17F52400";
    attribute INIT_16 of inst : label is "D555E1201B73A4E00959E6567BA90D49A6895521ABCA0268153D151F36AB93D9";
    attribute INIT_17 of inst : label is "1EF8CCD4A430D4B7B34333ED77ABF0466FFDFE7918C0F4001003315574CE9595";
    attribute INIT_18 of inst : label is "30343C1795C8552281054A0D55555E0142A40A303A9A0B05547E8294F6BFFA1F";
    attribute INIT_19 of inst : label is "F1FA5B6D54481A346563C0D0D5C55FF54A67F28FB96B32AB295C00158FA70B2B";
    attribute INIT_1A of inst : label is "0019A0D305916FC3D000400CC555D33A5657555784806DCE938025679959EEA5";
    attribute INIT_1B of inst : label is "63C2972FC140E0700B102508BD0FA600D62023ACFEC563F9C1CF0353CCC5729E";
    attribute INIT_1C of inst : label is "578AD958C574CC2EF89000009555425A0632B03FEAE80DD5575C014516355555";
    attribute INIT_1D of inst : label is "05C15728DAD082D3347B8F59A003C6B0557C47392E4AF8001B47FEF0A84AA785";
    attribute INIT_1E of inst : label is "4C5148000C1171B15555C39472C052B001BF0104FEFC0EBAC50F67ACC3FC3902";
    attribute INIT_1F of inst : label is "5AB2E502C5553A1BE8D012CF88001A5582C0C1FEBE3C018EC57A98FDF26A0542";
    attribute INIT_20 of inst : label is "0A8FA1275554CF21488003AFA6AFBC45575FBD80DB2F84A66FFE4A7D0357290A";
    attribute INIT_21 of inst : label is "C00AA006C06FFE5D5602AC555555C50C6A4C000B30F95BCEB1060D3D59635EED";
    attribute INIT_22 of inst : label is "0002AB6FB9F37E0C07C89ABDF333B340A444D021D5780000DFDB5241682AFEFD";
    attribute INIT_23 of inst : label is "1FFF3EC55736CF35EAAAFF9036BF8FB3FEEEF8F86C5955A1B15780664FF11A75";
    attribute INIT_24 of inst : label is "0444C093D952BACC550EA3EBB1012643300C7D5421500F50B4045028488179E6";
    attribute INIT_25 of inst : label is "C1A5540684AFF93806C300CF1BCF9A6816F0BBA54A97ECCEF1F555F912F9366D";
    attribute INIT_26 of inst : label is "FC2FFD6694E6AC930CF0A55270143102B28C96ABADAF95254CC0A64EA9AFC01F";
    attribute INIT_27 of inst : label is "990CC032F55784444A86214972A52E0129E56C333EC5830BFF83EBAC32500BBB";
    attribute INIT_28 of inst : label is "2A54498A3EE03A2BEACF161550E44BE4D9B41113024F654AEB31543A8FAEC404";
    attribute INIT_29 of inst : label is "B06F55EA84EAC3CD330EEF0BA3FBB6AEB103E1455C2FBEFE8290E8640CFBED3D";
    attribute INIT_2A of inst : label is "182B04F55873AEEBFDA90A6C46A90E669ECC57FF870C990EBFC395107548FFD9";
    attribute INIT_2B of inst : label is "D6BA40D33AECF006B37E849F147CE9816F07CFAA830EAD005F0CA43333CE4CC4";
    attribute INIT_2C of inst : label is "53E96E6800AAAAA6661EABBBF4FA6BAB311F8ED6BC1573E69A600F3BE83AA3FF";
    attribute INIT_2D of inst : label is "1A96000EA41C9A51CEAF2940510990401693EB565840FAEB53CC550454473282";
    attribute INIT_2E of inst : label is "C4AA5BE6A950EBE1669050C35BA90FC2440A8D9105047F000AFD4CE06AEB0511";
    attribute INIT_2F of inst : label is "BF5BBEA93F15A7EA9983C0FBAF05999507335A00CF38C0F1190010413FA6C03B";
    attribute INIT_30 of inst : label is "1443969BA6B30AFA9615530057FEF8CBF0143002F000033C30FF3459A800100C";
    attribute INIT_31 of inst : label is "40A045028101003BAFF35404544A6AA00CFEF303C4146A832ABCCF5AFB69943C";
    attribute INIT_32 of inst : label is "01104101511153FA0C33F041A9413FFCC0466910457CCC4573A8F0CCC3C0D451";
    attribute INIT_33 of inst : label is "113C0543F01C00011155170300335445510501010545F430C033F4140010FC30";
    attribute INIT_34 of inst : label is "6545FC3B0D53F000181C3CF1302699014F55153FBE83ABCF1459541430CC4699";
    attribute INIT_35 of inst : label is "FFF30119A44115F33115CEA3C333CF0304554444044514315CEABC3451051546";
    attribute INIT_36 of inst : label is "3F1540001550154013033C0C5004051CF0CC0451400544454FE830CFC106A504";
    attribute INIT_37 of inst : label is "3FC0C51513F001000FC030419441FF3C500D5045413F4104F01400404030C300";
    attribute INIT_38 of inst : label is "050C554000D111540CFCCCF5414015403C0404100430501FFC0CFF34542A5151";
    attribute INIT_39 of inst : label is "5010004CC545557F011540CF3F3FC1450555543FCC5050F3FC3100510114110F";
    attribute INIT_3A of inst : label is "0554000050555400044510004555CF3FF010000011540014505540053C3D4000";
    attribute INIT_3B of inst : label is "000D540005000C55055544155000000004000101555540015044101044000100";
    attribute INIT_3C of inst : label is "405503F0015454055400FFD550FC00011455000000C5554000001110C0554010";
    attribute INIT_3D of inst : label is "555540010040003F0054550055440311501140111543FFCFF000040001544004";
    attribute INIT_3E of inst : label is "000003C100005501570C300154050000411005101543F015554CC5557C515551";
    attribute INIT_3F of inst : label is "000C40111554555000050004100001555400FC01410100054400445000010454";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "22B347BFFEE8BB96A0897222A8A0E02A9DD0AEBC8B4FE536856AB7BA62B40825";
    attribute INIT_01 of inst : label is "FC8263B1AF000DBFF67FFC3BC14B00042E09F68A3B9A71946C8EA898A880C9C7";
    attribute INIT_02 of inst : label is "3F001013C10BFFFFEB05C35B8C98D86A8FF7C7F5CCC000E1FFFA400020F014FF";
    attribute INIT_03 of inst : label is "CEC5519A99BA80FC0002AAAA802280802895CB7FFFB5E0097DD94662ABDD51D6";
    attribute INIT_04 of inst : label is "C8A580039FFFF32397C0117D4217FF79000C76FDB2FFC2CCEA1A9FC15503FFFF";
    attribute INIT_05 of inst : label is "1FFD33A04C66A82B79FB5E13661501AFF0F1005681003DFFFFEA833AD5539E0C";
    attribute INIT_06 of inst : label is "AE5D4AAA99543EAA6A100902B866AE88E2801C3C000F00033F02009AAB07E08F";
    attribute INIT_07 of inst : label is "AFFFF774945EF9274DCCB81648C47EA4B9A79080C5315008FA8B8CD68AFFEEAA";
    attribute INIT_08 of inst : label is "026D017FFFDEAD5620ED393501FCEC2EFFFF0D4171D2C14324428AEBFC74001F";
    attribute INIT_09 of inst : label is "8B7F502DD600000859C218FFFDCB5F46802ABBFFFAA80AA0003155DBA2238001";
    attribute INIT_0A of inst : label is "AE0482BA2FA3C9801B70E8A009C6A029C88288240D5392AE69683437FC01CC91";
    attribute INIT_0B of inst : label is "33A2E9F52BDE4C200F7332F98D90A81F0F8643AFDD826CA09477EDCE0B7F2194";
    attribute INIT_0C of inst : label is "7D1A00AAEFFFEAA02A8000C5576E888E000409B405FFFF72FF5D83A429E40B32";
    attribute INIT_0D of inst : label is "AAAAA20BE8208408DC051E0A2B7FFCBD3757737F8CCFC900005EF80767FFF7AD";
    attribute INIT_0E of inst : label is "2A000AD80AE55DE9A3AC8F000349DFFC8D824463E624FFE089F9A85C002AAAAA";
    attribute INIT_0F of inst : label is "C0FFF983A1915A708070EAAA6644F3A9AAAA4C1D13CB08B5A6A02C2800008A80";
    attribute INIT_10 of inst : label is "007C3BE4403FDFF280C7D3E0D00003801DF03BFFFFF7DE4DE35C2B3A3800B70B";
    attribute INIT_11 of inst : label is "9740B80286CD2B5FF7FBDDCB5F10A4048B014FFFDF5A255FFD1FF57AAB91CEC0";
    attribute INIT_12 of inst : label is "729FDE3F01FA7F49800837F42F69F00DDEAB900C26F79A83FDC1804EB0DC6DB6";
    attribute INIT_13 of inst : label is "F0BEBDD82FFF9DEFD22400147E861F143F76905ABFFFD75EB300005A0B52FF91";
    attribute INIT_14 of inst : label is "FF7EB77B02BBC68E638AA5FFCFAF7D3E9D65816A8F051FFFC028EFDE387D3B10";
    attribute INIT_15 of inst : label is "B1255FB420C85C5E22AA21FFF20C000182A2455645062CC57EA3F0FF43DDB9FF";
    attribute INIT_16 of inst : label is "B0004997E4DDA6375FF39B81512183C6FBEA0042FEA7573EE0F5BD320E89B026";
    attribute INIT_17 of inst : label is "6C2EA8BEAE8229E51F40880694DEA846CFD4DCEEE60A897F6FFE94001C236AE2";
    attribute INIT_18 of inst : label is "577CA29E60A10049565A1D2400000CA1C97177A02F6F7C2F7E616A9E294A87B7";
    attribute INIT_19 of inst : label is "0385ACE401E56F81381155F8372777F7C53228372E3C815403D8029720F3FC89";
    attribute INIT_1A of inst : label is "0A1B2FCD7F4C98AA25FDBFFA5000708DAB8AC001265F937698DD7FCE6E054487";
    attribute INIT_1B of inst : label is "282A34B00148379FF492852E37087902A98548F28B8DE2A67C0557D02050394B";
    attribute INIT_1C of inst : label is "03A72C84F01C3758FAEFFFFDF0001C77DB834A08171F5B40036FFEB061900000";
    attribute INIT_1D of inst : label is "855409BD6F3ACA65D6F380ACF7FD0E3D0016EFD9931D0DFFCC6F7C0A224D5A10";
    attribute INIT_1E of inst : label is "48734DFFF76E291C00024263AAFD0C07FEC2A1A623AA03CD2728BA0548220C7F";
    attribute INIT_1F of inst : label is "87C847A25000F0994A0FC87D07FF65AAD580A354B42AAB238FF8B2082AE0D01E";
    attribute INIT_20 of inst : label is "780AF38D2803608E1AFFFF787B78CAD0015AC2DFE405AEF1C5FC6848FDBFC3AD";
    attribute INIT_21 of inst : label is "9FD775592ACD5CD20B2A850000006852E2617FF4AA042E23C98C7F035BC2A32C";
    attribute INIT_22 of inst : label is "FFF5DEE73BDD1400ADF2ED43200A6917A4662F73C03A7FFFE01306CB68BFA0DF";
    attribute INIT_23 of inst : label is "E8282BA5DE8477DF355528CFD34A62CBD4EE58059A7B77291C0328CEC009BAC8";
    attribute INIT_24 of inst : label is "2ECE8218A6A74F2D02740A3EC389399FDFD2DC01C3DA88074F53F89D34B4131B";
    attribute INIT_25 of inst : label is "21A754A40C07590DF1200A8219F5BFBD49823B85EFC092A389D000D3BA718333";
    attribute INIT_26 of inst : label is "2AA7556EB439F2102028082CC8BC8B8A1E0A635ED10DBF8FC02A2C61F6F0A23A";
    attribute INIT_27 of inst : label is "E67F7F4A700B0E66EFD984316BD8FADCC11AB8A823A5A8A357A2B6FA018F5E64";
    attribute INIT_28 of inst : label is "17039EC2746A2F569FA0B6400F4EE9C60CCCBB3A08629A9D3CB409D028FB0E24";
    attribute INIT_29 of inst : label is "6A6D0040269789F780A1102308A443FBE38ABB6550AF96762B4FF664A8A60C5D";
    attribute INIT_2A of inst : label is "468BD17552E0D3097F01AF18E42109916320D5FD2C023B83400ACAE8D0128824";
    attribute INIT_2B of inst : label is "9E1060300DBAA804151E0EE03E4A1EF4B20FF78800AB79AAFDD78C800A2B1751";
    attribute INIT_2C of inst : label is "D8B691962A2A002CCCB3FECC0CADB476BCC723A1C017FD6C10CAA88162AFF828";
    attribute INIT_2D of inst : label is "B8B4AAABF162BAD909F22348F923B84A9E189C7ED24A0F1EF208DDA6FE4C8014";
    attribute INIT_2E of inst : label is "2E00D9CC01D0B69B4C985000F12B0208E425E319A52CE20A2AFF629517BCADB3";
    attribute INIT_2F of inst : label is "E0F1B409223F84954E48228EF207BB1D8E2850A000AE2AA3B1AA3861A871208C";
    attribute INIT_30 of inst : label is "164AEB44D9C0A87A3CBFF0225D5450268ABE82AB820A22A28A2AA47BA282B82A";
    attribute INIT_31 of inst : label is "EA0A6F882303A88C5088D40E5C62428228210A000C1660AA9F6028D271C99E22";
    attribute INIT_32 of inst : label is "23B06B03F9BBF8AF20A028E10163A20AA2ECE390E5C8A06DC2FE802A000034F9";
    attribute INIT_33 of inst : label is "BB00256002B2A881B3D5BC82AAA8FCE55905A901A56F0C002AA28E3EA8B2A880";
    attribute INIT_34 of inst : label is "EF4708AE83F000089238AA83028EB1AB40F7B7A843EAD4881679F616080864B1";
    attribute INIT_35 of inst : label is "882A8BB38E43972281B70BFA00A8000024F7EE6EAE659C03F23FEA0E510F9564";
    attribute INIT_36 of inst : label is "809542A815703FC030AA80A2D2A6ADB2A2008ED1680FE6EFE2BC8280A384058E";
    attribute INIT_37 of inst : label is "002A0797BA8089A220000AC916CB2020F003F8E56100C98C0216A26868AA80A2";
    attribute INIT_38 of inst : label is "0F00FFC000333B7CAA82220D43EA97C002AE269A8400D2B22A8A000E54807B73";
    attribute INIT_39 of inst : label is "703028C0254557C0033FCAA0808003E5057FFC000050580AAA8300FB039E1B00";
    attribute INIT_3A of inst : label is "AFFC0000FAFFFC000EEFBAA0E5FF00AA003A800039FC003E5057C00F08234AA8";
    attribute INIT_3B of inst : label is "00015400250002550FFFCC3FF00008000E8003ABFFFFC003F8EE9ABAEEA823AA";
    attribute INIT_3C of inst : label is "E8FF000003D456AFFC00003FF0000029967F000000255FC0000039B020FFC030";
    attribute INIT_3D of inst : label is "FFFFC003AAC0000000FE55AAFFCC00B95AB3C03BBFC000200000A6AAABFCC00E";
    attribute INIT_3E of inst : label is "000000030000FFABFC000003FEAF0000EBB00FBABFC0003FFFC00FFFC0F3FFF3";
    attribute INIT_3F of inst : label is "0000C03BBFFCFFF0000F000EB00003FFFC000003EBAB000FEC00EEF00003AEFC";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "F396045FFE23B1A9050E430B0006A939E57716AA5390005AAAAC5AFFE95AA54E";
    attribute INIT_01 of inst : label is "FD4EA8D62EC00A4FFEFFE37FF81200056C6BF6D0541DE6E5748E40FB21C75171";
    attribute INIT_02 of inst : label is "71001ABADD7BFFFFED4D967EA6B2D48A1FFD1FFD1C4000E77FF0C00004389E7F";
    attribute INIT_03 of inst : label is "BABFFFFFFFFFC0FC0000000015441515553AD8FFFE5F2159FD6E5B04FE557EF9";
    attribute INIT_04 of inst : label is "16A80002BFFFF678FF2F60AB226AFFD000015B14C6FFD5FBDDF6002FFFFEAAAA";
    attribute INIT_05 of inst : label is "E69545D3669D541AA1156DA9AC8BB2BEC054001DC9000BFFFFA49CD07BFEA551";
    attribute INIT_06 of inst : label is "0E277FFFFFFFEAAAAAF1BF9CCBFFFFFBF0153BFC000F00033F005535AAFFC547";
    attribute INIT_07 of inst : label is "2DFFF838256D5543FABED29526BDFB2A42FEAAB19BAC90016213F3B048BFE200";
    attribute INIT_08 of inst : label is "E19EB2FFFF49DE5BB0FFEA95556D5EAD2FFFA655AC715B554D39BCD81BB40019";
    attribute INIT_09 of inst : label is "FFEAC8B2F0C0001C298725FFFE88E5DC1555555555555005551D6AB1C051D000";
    attribute INIT_0A of inst : label is "0EAB9558BFFD6A340EA16C003ABF1B03A51550EC0FFEA956C6903C8FFE5A7DFF";
    attribute INIT_0B of inst : label is "79B76BFDAE6B17052EAD6396BF7ABF7416DDB1ABE0E64C06BE2401879AFE13AC";
    attribute INIT_0C of inst : label is "977055555555555540155475AAC701474003867ACBFFFD27796EC3FFEA5555F5";
    attribute INIT_0D of inst : label is "0000045555050FFA515B6F9032BFFABF32AAAE96EEDBD200003CA71F97FFFA23";
    attribute INIT_0E of inst : label is "4000016A40C99E6A97446F00012E7FFE590071637F2AFF87BF96F92C00000000";
    attribute INIT_0F of inst : label is "AAFFC1FF7853F6ED83A0FFFFFFFFAEAAAAAAA00C0586E01B02296C0155555555";
    attribute INIT_10 of inst : label is "00222BEF800FFFFA06EFE1E9E00005DDF7C043FFFFFFF6C905ABF1FE47149101";
    attribute INIT_11 of inst : label is "A9555B1DA1E7552FEF31A0437544DAAB810153FFFA3DD2FFFFF55AD18B93D1C0";
    attribute INIT_12 of inst : label is "122FFAD64EFAFF5100137BFE414BD01659D9C4051B0B4F57FEE73C869DADEA2D";
    attribute INIT_13 of inst : label is "94FE28771FFF76CDF1640029B153ECE413BD31107FFFEAE18D00009A9ED5FDB3";
    attribute INIT_14 of inst : label is "FF896FD3F3929C17AB731E1561B54206AB8E012E5D0633FFB4072FE277AD9372";
    attribute INIT_15 of inst : label is "AE0ADDF95B1EF01861B95C7FF8BD00024395E2EC7947846BDE78816906C21EFF";
    attribute INIT_16 of inst : label is "54009B27E17B1B8AD60B7052CF0583DB0E7C00570E58A44A8012FAF04DFC12F3";
    attribute INIT_17 of inst : label is "0A15013A4215D988EB701518248E40F95EA569ED481571BFEFF58800131AFFC4";
    attribute INIT_18 of inst : label is "A9A304FD19B1004E1AAA936100001EAFC70A9D406C005225AACB896B1CE5BE61";
    attribute INIT_19 of inst : label is "032C3AC4025149617C2F41883F3E92B59B0292DB887506FE247153E462CA932E";
    attribute INIT_1A of inst : label is "53E57A51A3862015C6FFBFD620004C6BFF1150026C9F85EC6E2B582DC14B3C16";
    attribute INIT_1B of inst : label is "4C395C6F8FF8B5BFF1FEA614BCC1BE41B31839A9150F5C58FDB2062C54107E09";
    attribute INIT_1C of inst : label is "014AF29BD010DFC1A3AFFAFE440009B852459EC1BD62D58002FBFE5AA6F00000";
    attribute INIT_1D of inst : label is "39D0039EE13158818A7F7210C6FFC4D00012E2636C9EBDFFD4E25E1246D6CC50";
    attribute INIT_1E of inst : label is "80EFC6FFFDAA6384000036192C400497F754EFEB6EA55ABF65C6C1B637D319F6";
    attribute INIT_1F of inst : label is "CE491B0DC000769EB29BD6EB4EFF7C0F173C0CFFF20039A15D310B18DD198008";
    attribute INIT_20 of inst : label is "1DB297A2400035D8103FFE2BF026B8000776BF2F93606C72DFFDA58AFFF2B1DB";
    attribute INIT_21 of inst : label is "AFE2B693920F9724A2790D000001FE9C7C8DFFF2406D9D054AB744C3E422FD19";
    attribute INIT_22 of inst : label is "BFF7A5DEF0F95DD534A27F9305419B461BEB9FB590157FFF89365B43976AA1AE";
    attribute INIT_23 of inst : label is "4900054E6C5DE9775B0FD19BFBAA955B5BFC071D4881FD5A740285E0700F959E";
    attribute INIT_24 of inst : label is "FFBC0EADB157AABD005B18AA53FA1C1ABF9B49009FFA8719C106216D9C101D2C";
    attribute INIT_25 of inst : label is "9255ACE5BF93F223F8800014375B7701A3927F1BDB13A9555ED0018B39377012";
    attribute INIT_26 of inst : label is "40DDB1555B1CE7AC55537009D53D53F93B71B33AA77B1AA5814E41B6AF955431";
    attribute INIT_27 of inst : label is "706AFE6D24027FEADB27195DC5867191776CD00059396C27FF755A95462A9EAA";
    attribute INIT_28 of inst : label is "205A934B9B1B6C4EA55A7B40022CE4DDC04BFEF03AB6C55EAAF4016C62A94FE8";
    attribute INIT_29 of inst : label is "8E9E41B1AC6A98AC8506E927186AB39543C693EAB08AC3F061EF889BC1692919";
    attribute INIT_2A of inst : label is "9DE255B6AAC56D2EAC5A8849EA46C2C3FE95E4976C0381DAE4162A7725622BF0";
    attribute INIT_2B of inst : label is "3406C5306B95000E7958BDBE7AC1C01A2947AAC1B15593AA4E562BC5541B6FEA";
    attribute INIT_2C of inst : label is "2DAFFFF94E95555166B5556A4C183FFDB51B61B0F93E7AC6A9185648F62F95AA";
    attribute INIT_2D of inst : label is "8FC6BFC6CA77401B16A8D5BCFFE95BC0E56DB9D01AC1A5A4F05356AAAABC0DEB";
    attribute INIT_2E of inst : label is "4EAA50C156B15AA7916BF0149406154A6C5B92ABFFEBC43AE4FCB1854EAA4FF3";
    attribute INIT_2F of inst : label is "5494F156042418700F90056554394056BC40EAB0155555579AAAFFAF1BF39566";
    attribute INIT_30 of inst : label is "EAC1BF0FBFA4E53F06BFF054E0EBC71AA4EBC555543AF05400554F955ABEAC01";
    attribute INIT_31 of inst : label is "FEAAFFFAAF03FC16AA50FFFAABE9556F015AA4000FFE956C6A9555E430156C43";
    attribute INIT_32 of inst : label is "3EAFFF03FFFFF155400540FEAAAF05A503A505B0FFC100EBC555000000003FAB";
    attribute INIT_33 of inst : label is "AF003FF003F000FFF3FFFC140000FCFFFFFFFFFFFFFF0C0000040FEAABF00100";
    attribute INIT_34 of inst : label is "55BF015553F0000FAAF1550303A55AAAC0FEAF06A9556A503E955AFF0150EA5A";
    attribute INIT_35 of inst : label is "16940E9416C3FF0403AF1554000000003FAFFAABFFEABC03F055554FFFFABFEA";
    attribute INIT_36 of inst : label is "00FFFEABFFF03FC030000000FEAAABF00400FABFFC0FFFFFC555001503FAAABC";
    attribute INIT_37 of inst : label is "00000EAAF0150FF0555550FAAABF0540F003FFAAAF00FABC03FFFEABFC001554";
    attribute INIT_38 of inst : label is "0F00FFC00033EAFC0000000FFEAABFC0000FEAAABC00FFF05550000FFFA55AF3";
    attribute INIT_39 of inst : label is "F0303CC03FFFFFC0033FC000000003FFFFFFFC0000FFFC00000300FF03FAFF00";
    attribute INIT_3A of inst : label is "FFFC0000FFFFFC000FFFFFF0FFFF0000003FC0003FFC003FFFFFC00F0143FAAB";
    attribute INIT_3B of inst : label is "0003FC003F0003FF0FFFCC3FF0000C000FC003FFFFFFC003FCFFFFFFFFFC33FF";
    attribute INIT_3C of inst : label is "FCFF000003FFFFFFFC00003FF000003FFFFF0000003FFFC000003FF000FFC030";
    attribute INIT_3D of inst : label is "FFFFC003FFC0000000FFFFFFFFCC00FFFFF3C03FFFC000000000FFFFFFFCC00F";
    attribute INIT_3E of inst : label is "000000030000FFFFFC000003FFFF0000FFF00FFFFFC0003FFFC00FFFC0F3FFF3";
    attribute INIT_3F of inst : label is "0000C03FFFFCFFF0000F000FF00003FFFC000003FFFF000FFC00FFF00003FFFC";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "595401BFFFE95AAAAAA55455AAAAAA950005AAAAA95555555556AAAAAAAAAAA5";
    attribute INIT_01 of inst : label is "FFA55500550001BFFFFFFE9555540001ABFFFE555556A90006BAAA55AFA40005";
    attribute INIT_02 of inst : label is "940006FE5006FFFFFAA50055555ABFA5BFFFFFFFFA00001AFFFE00001BEA56FF";
    attribute INIT_03 of inst : label is "5555555555556A56AAAAAAAAAAAAAAAAAA956BFFFF905AABFF900055000006AA";
    attribute INIT_04 of inst : label is "555500006FFFFE95005540005AFFFFE4000000551BFFF90016A9555555555555";
    attribute INIT_05 of inst : label is "0000001AFFFAAAAAAFE4015556BFE95500000001640007FFFFFFA50005555555";
    attribute INIT_06 of inst : label is "A540555555555555555AAAA5155555555AAA9556AAA5AAA995AAAA9555556AA4";
    attribute INIT_07 of inst : label is "ABFFFFEA4001555400016FFFEAABFE955555555ABFE5000005A954056BFFFEAA";
    attribute INIT_08 of inst : label is "1AA55AFFFFFA50005A5555555556A556FFFFE400015AA4006BEAABA555400001";
    attribute INIT_09 of inst : label is "000016AFFE000002FFA45BFFFFA50016AAAAAAAAAAAAAAAAAA9000056AA90000";
    attribute INIT_0A of inst : label is "A5555556AAAAAA95500556AA9555AAFEAAAAAA56A55555556AAA96BFFFFFE500";
    attribute INIT_0B of inst : label is "955AFFFF900055AA9001AEAAAA9555400016AFFFFFA9515555400015BFFFE956";
    attribute INIT_0C of inst : label is "005AAAAAAAAAAAAAAAAAAA400015AAA400006A956BFFFFE9400169555555555A";
    attribute INIT_0D of inst : label is "AAAAAAAAAAAAA5555555AAAA9AFFFFFFD400000016BFF8000007FE906FFFFE94";
    attribute INIT_0E of inst : label is "AAAAAAAAAA6BFAAAA956A4000056FFFF90000559405BFFF955555556AAAAAAAA";
    attribute INIT_0F of inst : label is "1BFFF9005BFEA901695A55555555555555555551556AAAAAFE9556AAAAAAAAAA";
    attribute INIT_10 of inst : label is "0005AFF90001BFFEAABFFE5500000016A9001AFFFFFFFE500000055555AA5400";
    attribute INIT_11 of inst : label is "555555ABFE55AAFFF945556940016AAAA4006FFFF9416FFFFE40001ABFFEBE00";
    attribute INIT_12 of inst : label is "5AFFF9006BFFFFE40005AFFFFFF90000016A5001AAF9506FFFA9416AABFA5541";
    attribute INIT_13 of inst : label is "AA55415AFFFFEABA5A900006AFFEA50005AA9406FFFFFFFE50000015501BFF94";
    attribute INIT_14 of inst : label is "FFFAAAA9595416AAFE9456FFFE4000555550005550005FFFEAAAFFFE9401545A";
    attribute INIT_15 of inst : label is "AA9016AAAAFA40015AAAABFFFF90000069556FFA40006BFFFA9500000015ABFF";
    attribute INIT_16 of inst : label is "900015AFFE4055BFF955AFFE5055696AFA90001AFAABFFF90005555AA5015AAE";
    attribute INIT_17 of inst : label is "01AAAA9555AABFA5005AAA9006BAAA555000016BFAAAAFFFFFFE500005AAAABF";
    attribute INIT_18 of inst : label is "0005AA56FF940016FFFFFE94000001556AFFFAAAABFFFE95556AA555ABAAAA94";
    attribute INIT_19 of inst : label is "A9ABEA50006FFAAFEBE40016959554056AFEA9006BEAAAAA955AA9555ABFFE90";
    attribute INIT_1A of inst : label is "A955400005BFEAAABFFFFFF9400016AAAAFE400056BFF90156FFE556BFF94155";
    attribute INIT_1B of inst : label is "169556AAA556AFFFFE5555AA416AAAAAAE9006AAAAA556ABFF940056AA4006FA";
    attribute INIT_1C of inst : label is "006AAFF90006BFF905BFFFFF9000015BFEAAA56AAAAFF900006FFFFFFE400000";
    attribute INIT_1D of inst : label is "9500006BFE9AA50015405AFFBFFFA50000055405ABFAABFFFA5401A9556ABA40";
    attribute INIT_1E of inst : label is "6A556BFFFFFFE95000005AFFE500016FFEAA5555AAAAAAAA956ABE405AA9ABFE";
    attribute INIT_1F of inst : label is "BAA555A50000055005BFF9006BFFEBFAFE96A50005AA955AA54555ABA5550001";
    attribute INIT_20 of inst : label is "015AA95400005A5006FFFFEAAFEAAA40005AAAFFFE9556AE5001556BFF94056A";
    attribute INIT_21 of inst : label is "BFFEAFFEA950005BFE95500000001BFA416BFFFEAAABFAAAA5540169555AAA90";
    attribute INIT_22 of inst : label is "FFFEAA500500016A9505AAA9AAAAA4005555BFE90006FFFFFA94006955AAA901";
    attribute INIT_23 of inst : label is "FAAAAAA556A50005AAFAAABFFEAAAAA4000155ABFA55555540006A555AA5556B";
    attribute INIT_24 of inst : label is "5556A556AFFEAA90000056AAA955ABFFFFF9500015556AFFA4005AABFA4001AB";
    attribute INIT_25 of inst : label is "A9555655555405AFFFAAAAAA94005AFFFEA940556AFEAAAAA50000159545AFE9";
    attribute INIT_26 of inst : label is "AA50055555ABA956AAA940016A96A955405AAEEAA94055556AA5555AAAAAAA9A";
    attribute INIT_27 of inst : label is "AFFFFFE5400055556AFE90016ABFE90005ABAAAAAA955694005AAAAAAAFFFAAA";
    attribute INIT_28 of inst : label is "AFFFFEA40055ABFAAAAA940000565516BFA5555A955ABFFAAA4000015AAAA556";
    attribute INIT_29 of inst : label is "A550000556AAA5016AAAAA9456AAAEAAA96AA9555A5014055ABFFA556AAA9001";
    attribute INIT_2A of inst : label is "FA540005556AAA9001556BFA55556ABEAAAA550056A9556AAAAAFFE94005AAAF";
    attribute INIT_2B of inst : label is "95556A9AAAAAAAA5400156AA956ABFFFEAA400155AAAA9555000556AAAAAFFFF";
    attribute INIT_2C of inst : label is "56AAAAAAA5555555555AAAAAA6ABEAAA40005AAFAA9540155556AAA505AAAAAA";
    attribute INIT_2D of inst : label is "5015556ABFE95555AAAA55565555556A5556AA55556AAAAA5AA955555556A500";
    attribute INIT_2E of inst : label is "A5555515555AAAA955555AAA5555AAA556AAA95555556A9555015ABFFAAAA559";
    attribute INIT_2F of inst : label is "AA550555AA9556AFFAAAAAAAAA95555556AA555AAAAAAAA955555555AAAEAAAA";
    attribute INIT_30 of inst : label is "556AAAFAAAAA554055555AAA550015AAAA556AAAAA955AAAAAAAA555555556AA";
    attribute INIT_31 of inst : label is "5555555555A956AAAAAA555555555555AAAAAAAAA5555556AAAAAA55455556A9";
    attribute INIT_32 of inst : label is "955555A955555AAAAAAAAA555555AAAAA955555A556AAA556AAAAAAAAAAA9555";
    attribute INIT_33 of inst : label is "55AA955AA95AAA55595556AAAAAA5655555555555555A6AAAAAAA555555AAAAA";
    attribute INIT_34 of inst : label is "5555AAAAA95AAAA5555AAAA9A95555556A5555AAAAAAAAAA95555555AAAA5555";
    attribute INIT_35 of inst : label is "AAAAA555556955AAA955AAAAAAAAAAAA95555555555556A95AAAAAA555555555";
    attribute INIT_36 of inst : label is "AA555555555A956A9AAAAAAA5555555AAAAA555556A555556AAAAAAAA9555556";
    attribute INIT_37 of inst : label is "AAAAA5555AAAA55AAAAAAA555555AAAA5AA9555555AA5556A955555556AAAAAA";
    attribute INIT_38 of inst : label is "A5AA556AAA995556AAAAAAA55555556AAAA5555556AA555AAAAAAAA555555559";
    attribute INIT_39 of inst : label is "5A9A966A9555556AA9956AAAAAAAA955555556AAAA5556AAAAA9AA55A95555AA";
    attribute INIT_3A of inst : label is "5556AAAA555556AAA555555A5555AAAAAA956AAA9556AA9555556AA5AAA95555";
    attribute INIT_3B of inst : label is "AAA956AA95AAA955A55566955AAAA6AAA56AA95555556AA95655555555569955";
    attribute INIT_3C of inst : label is "5655AAAAA955555556AAAA955AAAAA955555AAAAAA95556AAAAA955AAA556A9A";
    attribute INIT_3D of inst : label is "55556AA9556AAAAAAA5555555566AA5555596A95556AAAAAAAAA555555566AA5";
    attribute INIT_3E of inst : label is "AAAAAAA9AAAA555556AAAAA95555AAAA555AA555556AAA95556AA5556A595559";
    attribute INIT_3F of inst : label is "AAAA6A955556555AAAA5AAA55AAAA95556AAAAA95555AAA556AA555AAAA95556";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
